
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"f0",x"fa",x"c2",x"87"),
    12 => (x"86",x"c0",x"c6",x"4e"),
    13 => (x"49",x"f0",x"fa",x"c2"),
    14 => (x"48",x"d0",x"e3",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"db",x"e3"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"4a",x"66",x"c4",x"1e"),
    47 => (x"51",x"12",x"48",x"71"),
    48 => (x"26",x"87",x"fb",x"05"),
    49 => (x"1e",x"73",x"1e",x"4f"),
    50 => (x"c0",x"02",x"9a",x"72"),
    51 => (x"48",x"c0",x"87",x"e7"),
    52 => (x"a9",x"72",x"4b",x"c1"),
    53 => (x"72",x"87",x"d1",x"06"),
    54 => (x"87",x"c9",x"06",x"82"),
    55 => (x"a9",x"72",x"83",x"73"),
    56 => (x"c3",x"87",x"f4",x"01"),
    57 => (x"3a",x"b2",x"c1",x"87"),
    58 => (x"89",x"03",x"a9",x"72"),
    59 => (x"c1",x"07",x"80",x"73"),
    60 => (x"f3",x"05",x"2b",x"2a"),
    61 => (x"26",x"4b",x"26",x"87"),
    62 => (x"1e",x"75",x"1e",x"4f"),
    63 => (x"b7",x"71",x"4d",x"c4"),
    64 => (x"b9",x"ff",x"04",x"a1"),
    65 => (x"bd",x"c3",x"81",x"c1"),
    66 => (x"a2",x"b7",x"72",x"07"),
    67 => (x"c1",x"ba",x"ff",x"04"),
    68 => (x"07",x"bd",x"c1",x"82"),
    69 => (x"c1",x"87",x"ee",x"fe"),
    70 => (x"b8",x"ff",x"04",x"2d"),
    71 => (x"2d",x"07",x"80",x"c1"),
    72 => (x"c1",x"b9",x"ff",x"04"),
    73 => (x"4d",x"26",x"07",x"81"),
    74 => (x"11",x"1e",x"4f",x"26"),
    75 => (x"08",x"d4",x"ff",x"48"),
    76 => (x"48",x"66",x"c4",x"78"),
    77 => (x"a6",x"c8",x"88",x"c1"),
    78 => (x"05",x"98",x"70",x"58"),
    79 => (x"4f",x"26",x"87",x"ed"),
    80 => (x"48",x"d4",x"ff",x"1e"),
    81 => (x"68",x"78",x"ff",x"c3"),
    82 => (x"48",x"66",x"c4",x"51"),
    83 => (x"a6",x"c8",x"88",x"c1"),
    84 => (x"05",x"98",x"70",x"58"),
    85 => (x"4f",x"26",x"87",x"eb"),
    86 => (x"ff",x"1e",x"73",x"1e"),
    87 => (x"ff",x"c3",x"4b",x"d4"),
    88 => (x"c3",x"4a",x"6b",x"7b"),
    89 => (x"49",x"6b",x"7b",x"ff"),
    90 => (x"b1",x"72",x"32",x"c8"),
    91 => (x"6b",x"7b",x"ff",x"c3"),
    92 => (x"71",x"31",x"c8",x"4a"),
    93 => (x"7b",x"ff",x"c3",x"b2"),
    94 => (x"32",x"c8",x"49",x"6b"),
    95 => (x"48",x"71",x"b1",x"72"),
    96 => (x"4d",x"26",x"87",x"c4"),
    97 => (x"4b",x"26",x"4c",x"26"),
    98 => (x"5e",x"0e",x"4f",x"26"),
    99 => (x"0e",x"5d",x"5c",x"5b"),
   100 => (x"d4",x"ff",x"4a",x"71"),
   101 => (x"c3",x"49",x"72",x"4c"),
   102 => (x"7c",x"71",x"99",x"ff"),
   103 => (x"bf",x"d0",x"e3",x"c2"),
   104 => (x"d0",x"87",x"c8",x"05"),
   105 => (x"30",x"c9",x"48",x"66"),
   106 => (x"d0",x"58",x"a6",x"d4"),
   107 => (x"29",x"d8",x"49",x"66"),
   108 => (x"71",x"99",x"ff",x"c3"),
   109 => (x"49",x"66",x"d0",x"7c"),
   110 => (x"ff",x"c3",x"29",x"d0"),
   111 => (x"d0",x"7c",x"71",x"99"),
   112 => (x"29",x"c8",x"49",x"66"),
   113 => (x"71",x"99",x"ff",x"c3"),
   114 => (x"49",x"66",x"d0",x"7c"),
   115 => (x"71",x"99",x"ff",x"c3"),
   116 => (x"d0",x"49",x"72",x"7c"),
   117 => (x"99",x"ff",x"c3",x"29"),
   118 => (x"4b",x"6c",x"7c",x"71"),
   119 => (x"4d",x"ff",x"f0",x"c9"),
   120 => (x"05",x"ab",x"ff",x"c3"),
   121 => (x"ff",x"c3",x"87",x"d0"),
   122 => (x"c1",x"4b",x"6c",x"7c"),
   123 => (x"87",x"c6",x"02",x"8d"),
   124 => (x"02",x"ab",x"ff",x"c3"),
   125 => (x"48",x"73",x"87",x"f0"),
   126 => (x"1e",x"87",x"c7",x"fe"),
   127 => (x"d4",x"ff",x"49",x"c0"),
   128 => (x"78",x"ff",x"c3",x"48"),
   129 => (x"c8",x"c3",x"81",x"c1"),
   130 => (x"f1",x"04",x"a9",x"b7"),
   131 => (x"1e",x"4f",x"26",x"87"),
   132 => (x"87",x"e7",x"1e",x"73"),
   133 => (x"4b",x"df",x"f8",x"c4"),
   134 => (x"ff",x"c0",x"1e",x"c0"),
   135 => (x"49",x"f7",x"c1",x"f0"),
   136 => (x"c4",x"87",x"e7",x"fd"),
   137 => (x"05",x"a8",x"c1",x"86"),
   138 => (x"ff",x"87",x"ea",x"c0"),
   139 => (x"ff",x"c3",x"48",x"d4"),
   140 => (x"c0",x"c0",x"c1",x"78"),
   141 => (x"1e",x"c0",x"c0",x"c0"),
   142 => (x"c1",x"f0",x"e1",x"c0"),
   143 => (x"c9",x"fd",x"49",x"e9"),
   144 => (x"70",x"86",x"c4",x"87"),
   145 => (x"87",x"ca",x"05",x"98"),
   146 => (x"c3",x"48",x"d4",x"ff"),
   147 => (x"48",x"c1",x"78",x"ff"),
   148 => (x"e6",x"fe",x"87",x"cb"),
   149 => (x"05",x"8b",x"c1",x"87"),
   150 => (x"c0",x"87",x"fd",x"fe"),
   151 => (x"87",x"e6",x"fc",x"48"),
   152 => (x"ff",x"1e",x"73",x"1e"),
   153 => (x"ff",x"c3",x"48",x"d4"),
   154 => (x"c0",x"4b",x"d3",x"78"),
   155 => (x"f0",x"ff",x"c0",x"1e"),
   156 => (x"fc",x"49",x"c1",x"c1"),
   157 => (x"86",x"c4",x"87",x"d4"),
   158 => (x"ca",x"05",x"98",x"70"),
   159 => (x"48",x"d4",x"ff",x"87"),
   160 => (x"c1",x"78",x"ff",x"c3"),
   161 => (x"fd",x"87",x"cb",x"48"),
   162 => (x"8b",x"c1",x"87",x"f1"),
   163 => (x"87",x"db",x"ff",x"05"),
   164 => (x"f1",x"fb",x"48",x"c0"),
   165 => (x"5b",x"5e",x"0e",x"87"),
   166 => (x"d4",x"ff",x"0e",x"5c"),
   167 => (x"87",x"db",x"fd",x"4c"),
   168 => (x"c0",x"1e",x"ea",x"c6"),
   169 => (x"c8",x"c1",x"f0",x"e1"),
   170 => (x"87",x"de",x"fb",x"49"),
   171 => (x"a8",x"c1",x"86",x"c4"),
   172 => (x"fe",x"87",x"c8",x"02"),
   173 => (x"48",x"c0",x"87",x"ea"),
   174 => (x"fa",x"87",x"e2",x"c1"),
   175 => (x"49",x"70",x"87",x"da"),
   176 => (x"99",x"ff",x"ff",x"cf"),
   177 => (x"02",x"a9",x"ea",x"c6"),
   178 => (x"d3",x"fe",x"87",x"c8"),
   179 => (x"c1",x"48",x"c0",x"87"),
   180 => (x"ff",x"c3",x"87",x"cb"),
   181 => (x"4b",x"f1",x"c0",x"7c"),
   182 => (x"70",x"87",x"f4",x"fc"),
   183 => (x"eb",x"c0",x"02",x"98"),
   184 => (x"c0",x"1e",x"c0",x"87"),
   185 => (x"fa",x"c1",x"f0",x"ff"),
   186 => (x"87",x"de",x"fa",x"49"),
   187 => (x"98",x"70",x"86",x"c4"),
   188 => (x"c3",x"87",x"d9",x"05"),
   189 => (x"49",x"6c",x"7c",x"ff"),
   190 => (x"7c",x"7c",x"ff",x"c3"),
   191 => (x"c0",x"c1",x"7c",x"7c"),
   192 => (x"87",x"c4",x"02",x"99"),
   193 => (x"87",x"d5",x"48",x"c1"),
   194 => (x"87",x"d1",x"48",x"c0"),
   195 => (x"c4",x"05",x"ab",x"c2"),
   196 => (x"c8",x"48",x"c0",x"87"),
   197 => (x"05",x"8b",x"c1",x"87"),
   198 => (x"c0",x"87",x"fd",x"fe"),
   199 => (x"87",x"e4",x"f9",x"48"),
   200 => (x"c2",x"1e",x"73",x"1e"),
   201 => (x"c1",x"48",x"d0",x"e3"),
   202 => (x"ff",x"4b",x"c7",x"78"),
   203 => (x"78",x"c2",x"48",x"d0"),
   204 => (x"ff",x"87",x"c8",x"fb"),
   205 => (x"78",x"c3",x"48",x"d0"),
   206 => (x"e5",x"c0",x"1e",x"c0"),
   207 => (x"49",x"c0",x"c1",x"d0"),
   208 => (x"c4",x"87",x"c7",x"f9"),
   209 => (x"05",x"a8",x"c1",x"86"),
   210 => (x"c2",x"4b",x"87",x"c1"),
   211 => (x"87",x"c5",x"05",x"ab"),
   212 => (x"f9",x"c0",x"48",x"c0"),
   213 => (x"05",x"8b",x"c1",x"87"),
   214 => (x"fc",x"87",x"d0",x"ff"),
   215 => (x"e3",x"c2",x"87",x"f7"),
   216 => (x"98",x"70",x"58",x"d4"),
   217 => (x"c1",x"87",x"cd",x"05"),
   218 => (x"f0",x"ff",x"c0",x"1e"),
   219 => (x"f8",x"49",x"d0",x"c1"),
   220 => (x"86",x"c4",x"87",x"d8"),
   221 => (x"c3",x"48",x"d4",x"ff"),
   222 => (x"e0",x"c4",x"78",x"ff"),
   223 => (x"d8",x"e3",x"c2",x"87"),
   224 => (x"48",x"d0",x"ff",x"58"),
   225 => (x"d4",x"ff",x"78",x"c2"),
   226 => (x"78",x"ff",x"c3",x"48"),
   227 => (x"f5",x"f7",x"48",x"c1"),
   228 => (x"5b",x"5e",x"0e",x"87"),
   229 => (x"71",x"0e",x"5d",x"5c"),
   230 => (x"4d",x"ff",x"c3",x"4a"),
   231 => (x"75",x"4c",x"d4",x"ff"),
   232 => (x"48",x"d0",x"ff",x"7c"),
   233 => (x"75",x"78",x"c3",x"c4"),
   234 => (x"c0",x"1e",x"72",x"7c"),
   235 => (x"d8",x"c1",x"f0",x"ff"),
   236 => (x"87",x"d6",x"f7",x"49"),
   237 => (x"98",x"70",x"86",x"c4"),
   238 => (x"c0",x"87",x"c5",x"02"),
   239 => (x"87",x"f0",x"c0",x"48"),
   240 => (x"fe",x"c3",x"7c",x"75"),
   241 => (x"1e",x"c0",x"c8",x"7c"),
   242 => (x"f5",x"49",x"66",x"d4"),
   243 => (x"86",x"c4",x"87",x"dc"),
   244 => (x"7c",x"75",x"7c",x"75"),
   245 => (x"da",x"d8",x"7c",x"75"),
   246 => (x"7c",x"75",x"4b",x"e0"),
   247 => (x"05",x"99",x"49",x"6c"),
   248 => (x"8b",x"c1",x"87",x"c5"),
   249 => (x"75",x"87",x"f3",x"05"),
   250 => (x"48",x"d0",x"ff",x"7c"),
   251 => (x"48",x"c1",x"78",x"c2"),
   252 => (x"1e",x"87",x"cf",x"f6"),
   253 => (x"ff",x"4a",x"d4",x"ff"),
   254 => (x"d1",x"c4",x"48",x"d0"),
   255 => (x"7a",x"ff",x"c3",x"78"),
   256 => (x"f8",x"05",x"89",x"c1"),
   257 => (x"1e",x"4f",x"26",x"87"),
   258 => (x"4b",x"71",x"1e",x"73"),
   259 => (x"df",x"cd",x"ee",x"c5"),
   260 => (x"48",x"d4",x"ff",x"4a"),
   261 => (x"68",x"78",x"ff",x"c3"),
   262 => (x"a8",x"fe",x"c3",x"48"),
   263 => (x"c1",x"87",x"c5",x"02"),
   264 => (x"87",x"ed",x"05",x"8a"),
   265 => (x"c5",x"05",x"9a",x"72"),
   266 => (x"c0",x"48",x"c0",x"87"),
   267 => (x"9b",x"73",x"87",x"ea"),
   268 => (x"c8",x"87",x"cc",x"02"),
   269 => (x"49",x"73",x"1e",x"66"),
   270 => (x"c4",x"87",x"c5",x"f4"),
   271 => (x"c8",x"87",x"c6",x"86"),
   272 => (x"ee",x"fe",x"49",x"66"),
   273 => (x"48",x"d4",x"ff",x"87"),
   274 => (x"78",x"78",x"ff",x"c3"),
   275 => (x"c5",x"05",x"9b",x"73"),
   276 => (x"48",x"d0",x"ff",x"87"),
   277 => (x"48",x"c1",x"78",x"d0"),
   278 => (x"1e",x"87",x"eb",x"f4"),
   279 => (x"4a",x"71",x"1e",x"73"),
   280 => (x"d4",x"ff",x"4b",x"c0"),
   281 => (x"78",x"ff",x"c3",x"48"),
   282 => (x"c4",x"48",x"d0",x"ff"),
   283 => (x"d4",x"ff",x"78",x"c3"),
   284 => (x"78",x"ff",x"c3",x"48"),
   285 => (x"ff",x"c0",x"1e",x"72"),
   286 => (x"49",x"d1",x"c1",x"f0"),
   287 => (x"c4",x"87",x"cb",x"f4"),
   288 => (x"05",x"98",x"70",x"86"),
   289 => (x"c0",x"c8",x"87",x"cd"),
   290 => (x"49",x"66",x"cc",x"1e"),
   291 => (x"c4",x"87",x"f8",x"fd"),
   292 => (x"ff",x"4b",x"70",x"86"),
   293 => (x"78",x"c2",x"48",x"d0"),
   294 => (x"e9",x"f3",x"48",x"73"),
   295 => (x"5b",x"5e",x"0e",x"87"),
   296 => (x"c0",x"0e",x"5d",x"5c"),
   297 => (x"f0",x"ff",x"c0",x"1e"),
   298 => (x"f3",x"49",x"c9",x"c1"),
   299 => (x"1e",x"d2",x"87",x"dc"),
   300 => (x"49",x"d8",x"e3",x"c2"),
   301 => (x"c8",x"87",x"d0",x"fd"),
   302 => (x"c1",x"4c",x"c0",x"86"),
   303 => (x"ac",x"b7",x"d2",x"84"),
   304 => (x"c2",x"87",x"f8",x"04"),
   305 => (x"bf",x"97",x"d8",x"e3"),
   306 => (x"99",x"c0",x"c3",x"49"),
   307 => (x"05",x"a9",x"c0",x"c1"),
   308 => (x"c2",x"87",x"e7",x"c0"),
   309 => (x"bf",x"97",x"df",x"e3"),
   310 => (x"c2",x"31",x"d0",x"49"),
   311 => (x"bf",x"97",x"e0",x"e3"),
   312 => (x"72",x"32",x"c8",x"4a"),
   313 => (x"e1",x"e3",x"c2",x"b1"),
   314 => (x"b1",x"4a",x"bf",x"97"),
   315 => (x"ff",x"cf",x"4c",x"71"),
   316 => (x"c1",x"9c",x"ff",x"ff"),
   317 => (x"c1",x"34",x"ca",x"84"),
   318 => (x"e3",x"c2",x"87",x"e7"),
   319 => (x"49",x"bf",x"97",x"e1"),
   320 => (x"99",x"c6",x"31",x"c1"),
   321 => (x"97",x"e2",x"e3",x"c2"),
   322 => (x"b7",x"c7",x"4a",x"bf"),
   323 => (x"c2",x"b1",x"72",x"2a"),
   324 => (x"bf",x"97",x"dd",x"e3"),
   325 => (x"9d",x"cf",x"4d",x"4a"),
   326 => (x"97",x"de",x"e3",x"c2"),
   327 => (x"9a",x"c3",x"4a",x"bf"),
   328 => (x"e3",x"c2",x"32",x"ca"),
   329 => (x"4b",x"bf",x"97",x"df"),
   330 => (x"b2",x"73",x"33",x"c2"),
   331 => (x"97",x"e0",x"e3",x"c2"),
   332 => (x"c0",x"c3",x"4b",x"bf"),
   333 => (x"2b",x"b7",x"c6",x"9b"),
   334 => (x"81",x"c2",x"b2",x"73"),
   335 => (x"30",x"71",x"48",x"c1"),
   336 => (x"48",x"c1",x"49",x"70"),
   337 => (x"4d",x"70",x"30",x"75"),
   338 => (x"84",x"c1",x"4c",x"72"),
   339 => (x"c0",x"c8",x"94",x"71"),
   340 => (x"cc",x"06",x"ad",x"b7"),
   341 => (x"b7",x"34",x"c1",x"87"),
   342 => (x"b7",x"c0",x"c8",x"2d"),
   343 => (x"f4",x"ff",x"01",x"ad"),
   344 => (x"f0",x"48",x"74",x"87"),
   345 => (x"5e",x"0e",x"87",x"dc"),
   346 => (x"0e",x"5d",x"5c",x"5b"),
   347 => (x"eb",x"c2",x"86",x"f8"),
   348 => (x"78",x"c0",x"48",x"fe"),
   349 => (x"1e",x"f6",x"e3",x"c2"),
   350 => (x"de",x"fb",x"49",x"c0"),
   351 => (x"70",x"86",x"c4",x"87"),
   352 => (x"87",x"c5",x"05",x"98"),
   353 => (x"ce",x"c9",x"48",x"c0"),
   354 => (x"c1",x"4d",x"c0",x"87"),
   355 => (x"c1",x"fa",x"c0",x"7e"),
   356 => (x"e4",x"c2",x"49",x"bf"),
   357 => (x"c8",x"71",x"4a",x"ec"),
   358 => (x"87",x"ce",x"eb",x"4b"),
   359 => (x"c2",x"05",x"98",x"70"),
   360 => (x"c0",x"7e",x"c0",x"87"),
   361 => (x"49",x"bf",x"fd",x"f9"),
   362 => (x"4a",x"c8",x"e5",x"c2"),
   363 => (x"ea",x"4b",x"c8",x"71"),
   364 => (x"98",x"70",x"87",x"f8"),
   365 => (x"c0",x"87",x"c2",x"05"),
   366 => (x"c0",x"02",x"6e",x"7e"),
   367 => (x"ea",x"c2",x"87",x"fd"),
   368 => (x"c2",x"4d",x"bf",x"fc"),
   369 => (x"bf",x"9f",x"f4",x"eb"),
   370 => (x"d6",x"c5",x"48",x"7e"),
   371 => (x"c7",x"05",x"a8",x"ea"),
   372 => (x"fc",x"ea",x"c2",x"87"),
   373 => (x"87",x"ce",x"4d",x"bf"),
   374 => (x"e9",x"ca",x"48",x"6e"),
   375 => (x"c5",x"02",x"a8",x"d5"),
   376 => (x"c7",x"48",x"c0",x"87"),
   377 => (x"e3",x"c2",x"87",x"f1"),
   378 => (x"49",x"75",x"1e",x"f6"),
   379 => (x"c4",x"87",x"ec",x"f9"),
   380 => (x"05",x"98",x"70",x"86"),
   381 => (x"48",x"c0",x"87",x"c5"),
   382 => (x"c0",x"87",x"dc",x"c7"),
   383 => (x"49",x"bf",x"fd",x"f9"),
   384 => (x"4a",x"c8",x"e5",x"c2"),
   385 => (x"e9",x"4b",x"c8",x"71"),
   386 => (x"98",x"70",x"87",x"e0"),
   387 => (x"c2",x"87",x"c8",x"05"),
   388 => (x"c1",x"48",x"fe",x"eb"),
   389 => (x"c0",x"87",x"da",x"78"),
   390 => (x"49",x"bf",x"c1",x"fa"),
   391 => (x"4a",x"ec",x"e4",x"c2"),
   392 => (x"e9",x"4b",x"c8",x"71"),
   393 => (x"98",x"70",x"87",x"c4"),
   394 => (x"87",x"c5",x"c0",x"02"),
   395 => (x"e6",x"c6",x"48",x"c0"),
   396 => (x"f4",x"eb",x"c2",x"87"),
   397 => (x"c1",x"49",x"bf",x"97"),
   398 => (x"c0",x"05",x"a9",x"d5"),
   399 => (x"eb",x"c2",x"87",x"cd"),
   400 => (x"49",x"bf",x"97",x"f5"),
   401 => (x"02",x"a9",x"ea",x"c2"),
   402 => (x"c0",x"87",x"c5",x"c0"),
   403 => (x"87",x"c7",x"c6",x"48"),
   404 => (x"97",x"f6",x"e3",x"c2"),
   405 => (x"c3",x"48",x"7e",x"bf"),
   406 => (x"c0",x"02",x"a8",x"e9"),
   407 => (x"48",x"6e",x"87",x"ce"),
   408 => (x"02",x"a8",x"eb",x"c3"),
   409 => (x"c0",x"87",x"c5",x"c0"),
   410 => (x"87",x"eb",x"c5",x"48"),
   411 => (x"97",x"c1",x"e4",x"c2"),
   412 => (x"05",x"99",x"49",x"bf"),
   413 => (x"c2",x"87",x"cc",x"c0"),
   414 => (x"bf",x"97",x"c2",x"e4"),
   415 => (x"02",x"a9",x"c2",x"49"),
   416 => (x"c0",x"87",x"c5",x"c0"),
   417 => (x"87",x"cf",x"c5",x"48"),
   418 => (x"97",x"c3",x"e4",x"c2"),
   419 => (x"eb",x"c2",x"48",x"bf"),
   420 => (x"4c",x"70",x"58",x"fa"),
   421 => (x"c2",x"88",x"c1",x"48"),
   422 => (x"c2",x"58",x"fe",x"eb"),
   423 => (x"bf",x"97",x"c4",x"e4"),
   424 => (x"c2",x"81",x"75",x"49"),
   425 => (x"bf",x"97",x"c5",x"e4"),
   426 => (x"72",x"32",x"c8",x"4a"),
   427 => (x"f0",x"c2",x"7e",x"a1"),
   428 => (x"78",x"6e",x"48",x"cb"),
   429 => (x"97",x"c6",x"e4",x"c2"),
   430 => (x"a6",x"c8",x"48",x"bf"),
   431 => (x"fe",x"eb",x"c2",x"58"),
   432 => (x"d4",x"c2",x"02",x"bf"),
   433 => (x"fd",x"f9",x"c0",x"87"),
   434 => (x"e5",x"c2",x"49",x"bf"),
   435 => (x"c8",x"71",x"4a",x"c8"),
   436 => (x"87",x"d6",x"e6",x"4b"),
   437 => (x"c0",x"02",x"98",x"70"),
   438 => (x"48",x"c0",x"87",x"c5"),
   439 => (x"c2",x"87",x"f8",x"c3"),
   440 => (x"4c",x"bf",x"f6",x"eb"),
   441 => (x"5c",x"df",x"f0",x"c2"),
   442 => (x"97",x"db",x"e4",x"c2"),
   443 => (x"31",x"c8",x"49",x"bf"),
   444 => (x"97",x"da",x"e4",x"c2"),
   445 => (x"49",x"a1",x"4a",x"bf"),
   446 => (x"97",x"dc",x"e4",x"c2"),
   447 => (x"32",x"d0",x"4a",x"bf"),
   448 => (x"c2",x"49",x"a1",x"72"),
   449 => (x"bf",x"97",x"dd",x"e4"),
   450 => (x"72",x"32",x"d8",x"4a"),
   451 => (x"66",x"c4",x"49",x"a1"),
   452 => (x"cb",x"f0",x"c2",x"91"),
   453 => (x"f0",x"c2",x"81",x"bf"),
   454 => (x"e4",x"c2",x"59",x"d3"),
   455 => (x"4a",x"bf",x"97",x"e3"),
   456 => (x"e4",x"c2",x"32",x"c8"),
   457 => (x"4b",x"bf",x"97",x"e2"),
   458 => (x"e4",x"c2",x"4a",x"a2"),
   459 => (x"4b",x"bf",x"97",x"e4"),
   460 => (x"a2",x"73",x"33",x"d0"),
   461 => (x"e5",x"e4",x"c2",x"4a"),
   462 => (x"cf",x"4b",x"bf",x"97"),
   463 => (x"73",x"33",x"d8",x"9b"),
   464 => (x"f0",x"c2",x"4a",x"a2"),
   465 => (x"f0",x"c2",x"5a",x"d7"),
   466 => (x"c2",x"4a",x"bf",x"d3"),
   467 => (x"c2",x"92",x"74",x"8a"),
   468 => (x"72",x"48",x"d7",x"f0"),
   469 => (x"ca",x"c1",x"78",x"a1"),
   470 => (x"c8",x"e4",x"c2",x"87"),
   471 => (x"c8",x"49",x"bf",x"97"),
   472 => (x"c7",x"e4",x"c2",x"31"),
   473 => (x"a1",x"4a",x"bf",x"97"),
   474 => (x"c6",x"ec",x"c2",x"49"),
   475 => (x"c2",x"ec",x"c2",x"59"),
   476 => (x"31",x"c5",x"49",x"bf"),
   477 => (x"c9",x"81",x"ff",x"c7"),
   478 => (x"df",x"f0",x"c2",x"29"),
   479 => (x"cd",x"e4",x"c2",x"59"),
   480 => (x"c8",x"4a",x"bf",x"97"),
   481 => (x"cc",x"e4",x"c2",x"32"),
   482 => (x"a2",x"4b",x"bf",x"97"),
   483 => (x"92",x"66",x"c4",x"4a"),
   484 => (x"f0",x"c2",x"82",x"6e"),
   485 => (x"f0",x"c2",x"5a",x"db"),
   486 => (x"78",x"c0",x"48",x"d3"),
   487 => (x"48",x"cf",x"f0",x"c2"),
   488 => (x"c2",x"78",x"a1",x"72"),
   489 => (x"c2",x"48",x"df",x"f0"),
   490 => (x"78",x"bf",x"d3",x"f0"),
   491 => (x"48",x"e3",x"f0",x"c2"),
   492 => (x"bf",x"d7",x"f0",x"c2"),
   493 => (x"fe",x"eb",x"c2",x"78"),
   494 => (x"c9",x"c0",x"02",x"bf"),
   495 => (x"c4",x"48",x"74",x"87"),
   496 => (x"c0",x"7e",x"70",x"30"),
   497 => (x"f0",x"c2",x"87",x"c9"),
   498 => (x"c4",x"48",x"bf",x"db"),
   499 => (x"c2",x"7e",x"70",x"30"),
   500 => (x"6e",x"48",x"c2",x"ec"),
   501 => (x"f8",x"48",x"c1",x"78"),
   502 => (x"26",x"4d",x"26",x"8e"),
   503 => (x"26",x"4b",x"26",x"4c"),
   504 => (x"5b",x"5e",x"0e",x"4f"),
   505 => (x"71",x"0e",x"5d",x"5c"),
   506 => (x"fe",x"eb",x"c2",x"4a"),
   507 => (x"87",x"cb",x"02",x"bf"),
   508 => (x"2b",x"c7",x"4b",x"72"),
   509 => (x"ff",x"c1",x"4c",x"72"),
   510 => (x"72",x"87",x"c9",x"9c"),
   511 => (x"72",x"2b",x"c8",x"4b"),
   512 => (x"9c",x"ff",x"c3",x"4c"),
   513 => (x"bf",x"cb",x"f0",x"c2"),
   514 => (x"f9",x"f9",x"c0",x"83"),
   515 => (x"d9",x"02",x"ab",x"bf"),
   516 => (x"fd",x"f9",x"c0",x"87"),
   517 => (x"f6",x"e3",x"c2",x"5b"),
   518 => (x"f0",x"49",x"73",x"1e"),
   519 => (x"86",x"c4",x"87",x"fd"),
   520 => (x"c5",x"05",x"98",x"70"),
   521 => (x"c0",x"48",x"c0",x"87"),
   522 => (x"eb",x"c2",x"87",x"e6"),
   523 => (x"d2",x"02",x"bf",x"fe"),
   524 => (x"c4",x"49",x"74",x"87"),
   525 => (x"f6",x"e3",x"c2",x"91"),
   526 => (x"cf",x"4d",x"69",x"81"),
   527 => (x"ff",x"ff",x"ff",x"ff"),
   528 => (x"74",x"87",x"cb",x"9d"),
   529 => (x"c2",x"91",x"c2",x"49"),
   530 => (x"9f",x"81",x"f6",x"e3"),
   531 => (x"48",x"75",x"4d",x"69"),
   532 => (x"0e",x"87",x"c6",x"fe"),
   533 => (x"5d",x"5c",x"5b",x"5e"),
   534 => (x"4d",x"71",x"1e",x"0e"),
   535 => (x"49",x"c1",x"1e",x"c0"),
   536 => (x"c4",x"87",x"fe",x"d0"),
   537 => (x"9c",x"4c",x"70",x"86"),
   538 => (x"87",x"c2",x"c1",x"02"),
   539 => (x"4a",x"c6",x"ec",x"c2"),
   540 => (x"df",x"ff",x"49",x"75"),
   541 => (x"98",x"70",x"87",x"d9"),
   542 => (x"87",x"f2",x"c0",x"02"),
   543 => (x"49",x"75",x"4a",x"74"),
   544 => (x"df",x"ff",x"4b",x"cb"),
   545 => (x"98",x"70",x"87",x"fe"),
   546 => (x"87",x"e2",x"c0",x"02"),
   547 => (x"9c",x"74",x"1e",x"c0"),
   548 => (x"c4",x"87",x"c7",x"02"),
   549 => (x"78",x"c0",x"48",x"a6"),
   550 => (x"a6",x"c4",x"87",x"c5"),
   551 => (x"c4",x"78",x"c1",x"48"),
   552 => (x"fc",x"cf",x"49",x"66"),
   553 => (x"70",x"86",x"c4",x"87"),
   554 => (x"fe",x"05",x"9c",x"4c"),
   555 => (x"48",x"74",x"87",x"fe"),
   556 => (x"87",x"e5",x"fc",x"26"),
   557 => (x"5c",x"5b",x"5e",x"0e"),
   558 => (x"86",x"f8",x"0e",x"5d"),
   559 => (x"05",x"9b",x"4b",x"71"),
   560 => (x"48",x"c0",x"87",x"c5"),
   561 => (x"c8",x"87",x"dd",x"c2"),
   562 => (x"7d",x"c0",x"4d",x"a3"),
   563 => (x"c7",x"02",x"66",x"d8"),
   564 => (x"97",x"66",x"d8",x"87"),
   565 => (x"87",x"c5",x"05",x"bf"),
   566 => (x"c7",x"c2",x"48",x"c0"),
   567 => (x"49",x"66",x"d8",x"87"),
   568 => (x"70",x"87",x"f0",x"fd"),
   569 => (x"c1",x"02",x"6e",x"7e"),
   570 => (x"49",x"6e",x"87",x"f8"),
   571 => (x"7d",x"69",x"81",x"dc"),
   572 => (x"81",x"da",x"49",x"6e"),
   573 => (x"9f",x"4c",x"a3",x"c4"),
   574 => (x"eb",x"c2",x"7c",x"69"),
   575 => (x"d0",x"02",x"bf",x"fe"),
   576 => (x"d4",x"49",x"6e",x"87"),
   577 => (x"49",x"69",x"9f",x"81"),
   578 => (x"ff",x"ff",x"c0",x"4a"),
   579 => (x"c2",x"32",x"d0",x"9a"),
   580 => (x"72",x"4a",x"c0",x"87"),
   581 => (x"80",x"6c",x"48",x"49"),
   582 => (x"7b",x"c0",x"7c",x"70"),
   583 => (x"6c",x"49",x"a3",x"cc"),
   584 => (x"49",x"a3",x"d0",x"79"),
   585 => (x"a6",x"c4",x"79",x"c0"),
   586 => (x"d4",x"78",x"c0",x"48"),
   587 => (x"66",x"c4",x"4a",x"a3"),
   588 => (x"72",x"91",x"c8",x"49"),
   589 => (x"41",x"c0",x"49",x"a1"),
   590 => (x"66",x"c4",x"79",x"6c"),
   591 => (x"c8",x"80",x"c1",x"48"),
   592 => (x"b7",x"c6",x"58",x"a6"),
   593 => (x"e2",x"ff",x"04",x"a8"),
   594 => (x"c9",x"4a",x"6d",x"87"),
   595 => (x"c0",x"49",x"72",x"2a"),
   596 => (x"dd",x"ff",x"4a",x"f0"),
   597 => (x"4a",x"70",x"87",x"ef"),
   598 => (x"49",x"a3",x"c4",x"c1"),
   599 => (x"48",x"6e",x"79",x"72"),
   600 => (x"48",x"c0",x"87",x"c2"),
   601 => (x"f0",x"f9",x"8e",x"f8"),
   602 => (x"5b",x"5e",x"0e",x"87"),
   603 => (x"71",x"0e",x"5d",x"5c"),
   604 => (x"f9",x"f9",x"c0",x"4c"),
   605 => (x"74",x"78",x"ff",x"48"),
   606 => (x"ca",x"c1",x"02",x"9c"),
   607 => (x"49",x"a4",x"c8",x"87"),
   608 => (x"c2",x"c1",x"02",x"69"),
   609 => (x"4a",x"66",x"d0",x"87"),
   610 => (x"d4",x"82",x"49",x"6c"),
   611 => (x"66",x"d0",x"5a",x"a6"),
   612 => (x"eb",x"c2",x"b9",x"4d"),
   613 => (x"ff",x"4a",x"bf",x"fa"),
   614 => (x"71",x"99",x"72",x"ba"),
   615 => (x"e4",x"c0",x"02",x"99"),
   616 => (x"4b",x"a4",x"c4",x"87"),
   617 => (x"f8",x"f8",x"49",x"6b"),
   618 => (x"c2",x"7b",x"70",x"87"),
   619 => (x"49",x"bf",x"f6",x"eb"),
   620 => (x"7c",x"71",x"81",x"6c"),
   621 => (x"eb",x"c2",x"b9",x"75"),
   622 => (x"ff",x"4a",x"bf",x"fa"),
   623 => (x"71",x"99",x"72",x"ba"),
   624 => (x"dc",x"ff",x"05",x"99"),
   625 => (x"f8",x"7c",x"75",x"87"),
   626 => (x"73",x"1e",x"87",x"cf"),
   627 => (x"9b",x"4b",x"71",x"1e"),
   628 => (x"c8",x"87",x"c7",x"02"),
   629 => (x"05",x"69",x"49",x"a3"),
   630 => (x"48",x"c0",x"87",x"c5"),
   631 => (x"c2",x"87",x"eb",x"c0"),
   632 => (x"4a",x"bf",x"cf",x"f0"),
   633 => (x"69",x"49",x"a3",x"c4"),
   634 => (x"c2",x"89",x"c2",x"49"),
   635 => (x"91",x"bf",x"f6",x"eb"),
   636 => (x"c2",x"4a",x"a2",x"71"),
   637 => (x"49",x"bf",x"fa",x"eb"),
   638 => (x"a2",x"71",x"99",x"6b"),
   639 => (x"1e",x"66",x"c8",x"4a"),
   640 => (x"d6",x"e9",x"49",x"72"),
   641 => (x"70",x"86",x"c4",x"87"),
   642 => (x"d0",x"f7",x"48",x"49"),
   643 => (x"1e",x"73",x"1e",x"87"),
   644 => (x"02",x"9b",x"4b",x"71"),
   645 => (x"a3",x"c8",x"87",x"c7"),
   646 => (x"c5",x"05",x"69",x"49"),
   647 => (x"c0",x"48",x"c0",x"87"),
   648 => (x"f0",x"c2",x"87",x"eb"),
   649 => (x"c4",x"4a",x"bf",x"cf"),
   650 => (x"49",x"69",x"49",x"a3"),
   651 => (x"eb",x"c2",x"89",x"c2"),
   652 => (x"71",x"91",x"bf",x"f6"),
   653 => (x"eb",x"c2",x"4a",x"a2"),
   654 => (x"6b",x"49",x"bf",x"fa"),
   655 => (x"4a",x"a2",x"71",x"99"),
   656 => (x"72",x"1e",x"66",x"c8"),
   657 => (x"87",x"c9",x"e5",x"49"),
   658 => (x"49",x"70",x"86",x"c4"),
   659 => (x"87",x"cd",x"f6",x"48"),
   660 => (x"5c",x"5b",x"5e",x"0e"),
   661 => (x"86",x"f8",x"0e",x"5d"),
   662 => (x"a6",x"c4",x"4b",x"71"),
   663 => (x"c8",x"78",x"ff",x"48"),
   664 => (x"4d",x"69",x"49",x"a3"),
   665 => (x"a3",x"d4",x"4c",x"c0"),
   666 => (x"c8",x"49",x"74",x"4a"),
   667 => (x"49",x"a1",x"72",x"91"),
   668 => (x"66",x"d8",x"49",x"69"),
   669 => (x"70",x"88",x"71",x"48"),
   670 => (x"a9",x"66",x"d8",x"7e"),
   671 => (x"6e",x"87",x"ca",x"01"),
   672 => (x"87",x"c5",x"06",x"ad"),
   673 => (x"6e",x"5c",x"a6",x"c8"),
   674 => (x"c6",x"84",x"c1",x"4d"),
   675 => (x"ff",x"04",x"ac",x"b7"),
   676 => (x"66",x"c4",x"87",x"d4"),
   677 => (x"f4",x"8e",x"f8",x"48"),
   678 => (x"5e",x"0e",x"87",x"ff"),
   679 => (x"0e",x"5d",x"5c",x"5b"),
   680 => (x"a6",x"c8",x"86",x"ec"),
   681 => (x"48",x"a6",x"c8",x"59"),
   682 => (x"ff",x"ff",x"ff",x"c1"),
   683 => (x"c4",x"78",x"ff",x"ff"),
   684 => (x"c0",x"78",x"ff",x"80"),
   685 => (x"c4",x"4c",x"c0",x"4d"),
   686 => (x"83",x"d4",x"4b",x"66"),
   687 => (x"91",x"c8",x"49",x"74"),
   688 => (x"75",x"49",x"a1",x"73"),
   689 => (x"73",x"92",x"c8",x"4a"),
   690 => (x"49",x"69",x"7e",x"a2"),
   691 => (x"d4",x"89",x"bf",x"6e"),
   692 => (x"ad",x"74",x"59",x"a6"),
   693 => (x"d0",x"87",x"c6",x"05"),
   694 => (x"bf",x"6e",x"48",x"a6"),
   695 => (x"48",x"66",x"d0",x"78"),
   696 => (x"04",x"a8",x"b7",x"c0"),
   697 => (x"66",x"d0",x"87",x"cf"),
   698 => (x"a9",x"66",x"c8",x"49"),
   699 => (x"d0",x"87",x"c6",x"03"),
   700 => (x"a6",x"cc",x"5c",x"a6"),
   701 => (x"c6",x"84",x"c1",x"59"),
   702 => (x"fe",x"04",x"ac",x"b7"),
   703 => (x"85",x"c1",x"87",x"f9"),
   704 => (x"04",x"ad",x"b7",x"c6"),
   705 => (x"cc",x"87",x"ee",x"fe"),
   706 => (x"8e",x"ec",x"48",x"66"),
   707 => (x"0e",x"87",x"ca",x"f3"),
   708 => (x"5d",x"5c",x"5b",x"5e"),
   709 => (x"71",x"86",x"f0",x"0e"),
   710 => (x"66",x"e0",x"c0",x"4b"),
   711 => (x"73",x"2c",x"c9",x"4c"),
   712 => (x"e1",x"c3",x"02",x"9b"),
   713 => (x"49",x"a3",x"c8",x"87"),
   714 => (x"d9",x"c3",x"02",x"69"),
   715 => (x"49",x"a3",x"d0",x"87"),
   716 => (x"79",x"66",x"e0",x"c0"),
   717 => (x"02",x"ac",x"7e",x"6b"),
   718 => (x"c2",x"87",x"cb",x"c3"),
   719 => (x"49",x"bf",x"fa",x"eb"),
   720 => (x"4a",x"71",x"b9",x"ff"),
   721 => (x"48",x"71",x"9a",x"74"),
   722 => (x"a6",x"cc",x"98",x"6e"),
   723 => (x"4d",x"a3",x"c4",x"58"),
   724 => (x"6d",x"48",x"a6",x"c4"),
   725 => (x"aa",x"66",x"c8",x"78"),
   726 => (x"74",x"87",x"c5",x"05"),
   727 => (x"87",x"d1",x"c2",x"7b"),
   728 => (x"49",x"73",x"1e",x"72"),
   729 => (x"c4",x"87",x"e9",x"fb"),
   730 => (x"48",x"7e",x"70",x"86"),
   731 => (x"04",x"a8",x"b7",x"c0"),
   732 => (x"a3",x"d4",x"87",x"d0"),
   733 => (x"c8",x"49",x"6e",x"4a"),
   734 => (x"49",x"a1",x"72",x"91"),
   735 => (x"7d",x"69",x"7b",x"21"),
   736 => (x"7b",x"c0",x"87",x"c7"),
   737 => (x"69",x"49",x"a3",x"cc"),
   738 => (x"1e",x"66",x"c8",x"7d"),
   739 => (x"ff",x"fa",x"49",x"73"),
   740 => (x"70",x"86",x"c4",x"87"),
   741 => (x"a3",x"c4",x"c1",x"7e"),
   742 => (x"48",x"a6",x"cc",x"49"),
   743 => (x"66",x"c8",x"78",x"69"),
   744 => (x"a8",x"66",x"cc",x"48"),
   745 => (x"6e",x"87",x"c9",x"06"),
   746 => (x"a8",x"b7",x"c0",x"48"),
   747 => (x"87",x"e0",x"c0",x"04"),
   748 => (x"b7",x"c0",x"48",x"6e"),
   749 => (x"ec",x"c0",x"04",x"a8"),
   750 => (x"4a",x"a3",x"d4",x"87"),
   751 => (x"91",x"c8",x"49",x"6e"),
   752 => (x"c8",x"49",x"a1",x"72"),
   753 => (x"88",x"69",x"48",x"66"),
   754 => (x"66",x"cc",x"49",x"70"),
   755 => (x"87",x"d5",x"06",x"a9"),
   756 => (x"c5",x"fb",x"49",x"73"),
   757 => (x"d4",x"49",x"70",x"87"),
   758 => (x"91",x"c8",x"4a",x"a3"),
   759 => (x"c8",x"49",x"a1",x"72"),
   760 => (x"66",x"c4",x"41",x"66"),
   761 => (x"74",x"8c",x"6b",x"79"),
   762 => (x"49",x"73",x"1e",x"49"),
   763 => (x"c4",x"87",x"fa",x"f5"),
   764 => (x"66",x"e0",x"c0",x"86"),
   765 => (x"99",x"ff",x"c7",x"49"),
   766 => (x"c2",x"87",x"cb",x"02"),
   767 => (x"73",x"1e",x"f6",x"e3"),
   768 => (x"87",x"c6",x"f7",x"49"),
   769 => (x"8e",x"f0",x"86",x"c4"),
   770 => (x"1e",x"87",x"ce",x"ef"),
   771 => (x"4b",x"71",x"1e",x"73"),
   772 => (x"e4",x"c0",x"02",x"9b"),
   773 => (x"e3",x"f0",x"c2",x"87"),
   774 => (x"c2",x"4a",x"73",x"5b"),
   775 => (x"f6",x"eb",x"c2",x"8a"),
   776 => (x"c2",x"92",x"49",x"bf"),
   777 => (x"48",x"bf",x"cf",x"f0"),
   778 => (x"f0",x"c2",x"80",x"72"),
   779 => (x"48",x"71",x"58",x"e7"),
   780 => (x"ec",x"c2",x"30",x"c4"),
   781 => (x"ed",x"c0",x"58",x"c6"),
   782 => (x"df",x"f0",x"c2",x"87"),
   783 => (x"d3",x"f0",x"c2",x"48"),
   784 => (x"f0",x"c2",x"78",x"bf"),
   785 => (x"f0",x"c2",x"48",x"e3"),
   786 => (x"c2",x"78",x"bf",x"d7"),
   787 => (x"02",x"bf",x"fe",x"eb"),
   788 => (x"eb",x"c2",x"87",x"c9"),
   789 => (x"c4",x"49",x"bf",x"f6"),
   790 => (x"c2",x"87",x"c7",x"31"),
   791 => (x"49",x"bf",x"db",x"f0"),
   792 => (x"ec",x"c2",x"31",x"c4"),
   793 => (x"f4",x"ed",x"59",x"c6"),
   794 => (x"5b",x"5e",x"0e",x"87"),
   795 => (x"4a",x"71",x"0e",x"5c"),
   796 => (x"9a",x"72",x"4b",x"c0"),
   797 => (x"87",x"e1",x"c0",x"02"),
   798 => (x"9f",x"49",x"a2",x"da"),
   799 => (x"eb",x"c2",x"4b",x"69"),
   800 => (x"cf",x"02",x"bf",x"fe"),
   801 => (x"49",x"a2",x"d4",x"87"),
   802 => (x"4c",x"49",x"69",x"9f"),
   803 => (x"9c",x"ff",x"ff",x"c0"),
   804 => (x"87",x"c2",x"34",x"d0"),
   805 => (x"49",x"74",x"4c",x"c0"),
   806 => (x"fd",x"49",x"73",x"b3"),
   807 => (x"fa",x"ec",x"87",x"ed"),
   808 => (x"5b",x"5e",x"0e",x"87"),
   809 => (x"f4",x"0e",x"5d",x"5c"),
   810 => (x"c0",x"4a",x"71",x"86"),
   811 => (x"02",x"9a",x"72",x"7e"),
   812 => (x"e3",x"c2",x"87",x"d8"),
   813 => (x"78",x"c0",x"48",x"f2"),
   814 => (x"48",x"ea",x"e3",x"c2"),
   815 => (x"bf",x"e3",x"f0",x"c2"),
   816 => (x"ee",x"e3",x"c2",x"78"),
   817 => (x"df",x"f0",x"c2",x"48"),
   818 => (x"ec",x"c2",x"78",x"bf"),
   819 => (x"50",x"c0",x"48",x"d3"),
   820 => (x"bf",x"c2",x"ec",x"c2"),
   821 => (x"f2",x"e3",x"c2",x"49"),
   822 => (x"aa",x"71",x"4a",x"bf"),
   823 => (x"87",x"c0",x"c4",x"03"),
   824 => (x"99",x"cf",x"49",x"72"),
   825 => (x"87",x"e1",x"c0",x"05"),
   826 => (x"1e",x"f6",x"e3",x"c2"),
   827 => (x"bf",x"ea",x"e3",x"c2"),
   828 => (x"ea",x"e3",x"c2",x"49"),
   829 => (x"78",x"a1",x"c1",x"48"),
   830 => (x"de",x"dd",x"ff",x"71"),
   831 => (x"c0",x"86",x"c4",x"87"),
   832 => (x"c2",x"48",x"f5",x"f9"),
   833 => (x"cc",x"78",x"f6",x"e3"),
   834 => (x"f5",x"f9",x"c0",x"87"),
   835 => (x"e0",x"c0",x"48",x"bf"),
   836 => (x"f9",x"f9",x"c0",x"80"),
   837 => (x"f2",x"e3",x"c2",x"58"),
   838 => (x"80",x"c1",x"48",x"bf"),
   839 => (x"58",x"f6",x"e3",x"c2"),
   840 => (x"00",x"0e",x"75",x"27"),
   841 => (x"bf",x"97",x"bf",x"00"),
   842 => (x"c2",x"02",x"9d",x"4d"),
   843 => (x"e5",x"c3",x"87",x"e2"),
   844 => (x"db",x"c2",x"02",x"ad"),
   845 => (x"f5",x"f9",x"c0",x"87"),
   846 => (x"a3",x"cb",x"4b",x"bf"),
   847 => (x"cf",x"4c",x"11",x"49"),
   848 => (x"d2",x"c1",x"05",x"ac"),
   849 => (x"df",x"49",x"75",x"87"),
   850 => (x"cd",x"89",x"c1",x"99"),
   851 => (x"c6",x"ec",x"c2",x"91"),
   852 => (x"4a",x"a3",x"c1",x"81"),
   853 => (x"a3",x"c3",x"51",x"12"),
   854 => (x"c5",x"51",x"12",x"4a"),
   855 => (x"51",x"12",x"4a",x"a3"),
   856 => (x"12",x"4a",x"a3",x"c7"),
   857 => (x"4a",x"a3",x"c9",x"51"),
   858 => (x"a3",x"ce",x"51",x"12"),
   859 => (x"d0",x"51",x"12",x"4a"),
   860 => (x"51",x"12",x"4a",x"a3"),
   861 => (x"12",x"4a",x"a3",x"d2"),
   862 => (x"4a",x"a3",x"d4",x"51"),
   863 => (x"a3",x"d6",x"51",x"12"),
   864 => (x"d8",x"51",x"12",x"4a"),
   865 => (x"51",x"12",x"4a",x"a3"),
   866 => (x"12",x"4a",x"a3",x"dc"),
   867 => (x"4a",x"a3",x"de",x"51"),
   868 => (x"7e",x"c1",x"51",x"12"),
   869 => (x"74",x"87",x"f9",x"c0"),
   870 => (x"05",x"99",x"c8",x"49"),
   871 => (x"74",x"87",x"ea",x"c0"),
   872 => (x"05",x"99",x"d0",x"49"),
   873 => (x"66",x"dc",x"87",x"d0"),
   874 => (x"87",x"ca",x"c0",x"02"),
   875 => (x"66",x"dc",x"49",x"73"),
   876 => (x"02",x"98",x"70",x"0f"),
   877 => (x"05",x"6e",x"87",x"d3"),
   878 => (x"c2",x"87",x"c6",x"c0"),
   879 => (x"c0",x"48",x"c6",x"ec"),
   880 => (x"f5",x"f9",x"c0",x"50"),
   881 => (x"e7",x"c2",x"48",x"bf"),
   882 => (x"d3",x"ec",x"c2",x"87"),
   883 => (x"7e",x"50",x"c0",x"48"),
   884 => (x"bf",x"c2",x"ec",x"c2"),
   885 => (x"f2",x"e3",x"c2",x"49"),
   886 => (x"aa",x"71",x"4a",x"bf"),
   887 => (x"87",x"c0",x"fc",x"04"),
   888 => (x"bf",x"e3",x"f0",x"c2"),
   889 => (x"87",x"c8",x"c0",x"05"),
   890 => (x"bf",x"fe",x"eb",x"c2"),
   891 => (x"87",x"fe",x"c1",x"02"),
   892 => (x"48",x"f9",x"f9",x"c0"),
   893 => (x"e3",x"c2",x"78",x"ff"),
   894 => (x"e7",x"49",x"bf",x"ee"),
   895 => (x"49",x"70",x"87",x"e3"),
   896 => (x"59",x"f2",x"e3",x"c2"),
   897 => (x"c2",x"48",x"a6",x"c4"),
   898 => (x"78",x"bf",x"ee",x"e3"),
   899 => (x"bf",x"fe",x"eb",x"c2"),
   900 => (x"87",x"d8",x"c0",x"02"),
   901 => (x"cf",x"49",x"66",x"c4"),
   902 => (x"f8",x"ff",x"ff",x"ff"),
   903 => (x"c0",x"02",x"a9",x"99"),
   904 => (x"4d",x"c0",x"87",x"c5"),
   905 => (x"c1",x"87",x"e1",x"c0"),
   906 => (x"87",x"dc",x"c0",x"4d"),
   907 => (x"cf",x"49",x"66",x"c4"),
   908 => (x"a9",x"99",x"f8",x"ff"),
   909 => (x"87",x"c8",x"c0",x"02"),
   910 => (x"c0",x"48",x"a6",x"c8"),
   911 => (x"87",x"c5",x"c0",x"78"),
   912 => (x"c1",x"48",x"a6",x"c8"),
   913 => (x"4d",x"66",x"c8",x"78"),
   914 => (x"c0",x"05",x"9d",x"75"),
   915 => (x"66",x"c4",x"87",x"e0"),
   916 => (x"c2",x"89",x"c2",x"49"),
   917 => (x"4a",x"bf",x"f6",x"eb"),
   918 => (x"cf",x"f0",x"c2",x"91"),
   919 => (x"e3",x"c2",x"4a",x"bf"),
   920 => (x"a1",x"72",x"48",x"ea"),
   921 => (x"f2",x"e3",x"c2",x"78"),
   922 => (x"f9",x"78",x"c0",x"48"),
   923 => (x"48",x"c0",x"87",x"e2"),
   924 => (x"e4",x"e5",x"8e",x"f4"),
   925 => (x"00",x"00",x"00",x"87"),
   926 => (x"ff",x"ff",x"ff",x"00"),
   927 => (x"00",x"0e",x"85",x"ff"),
   928 => (x"00",x"0e",x"8e",x"00"),
   929 => (x"54",x"41",x"46",x"00"),
   930 => (x"20",x"20",x"32",x"33"),
   931 => (x"41",x"46",x"00",x"20"),
   932 => (x"20",x"36",x"31",x"54"),
   933 => (x"1e",x"00",x"20",x"20"),
   934 => (x"c3",x"48",x"d4",x"ff"),
   935 => (x"48",x"68",x"78",x"ff"),
   936 => (x"ff",x"1e",x"4f",x"26"),
   937 => (x"ff",x"c3",x"48",x"d4"),
   938 => (x"48",x"d0",x"ff",x"78"),
   939 => (x"ff",x"78",x"e1",x"c8"),
   940 => (x"78",x"d4",x"48",x"d4"),
   941 => (x"48",x"e7",x"f0",x"c2"),
   942 => (x"50",x"bf",x"d4",x"ff"),
   943 => (x"ff",x"1e",x"4f",x"26"),
   944 => (x"e0",x"c0",x"48",x"d0"),
   945 => (x"1e",x"4f",x"26",x"78"),
   946 => (x"70",x"87",x"cc",x"ff"),
   947 => (x"c6",x"02",x"99",x"49"),
   948 => (x"a9",x"fb",x"c0",x"87"),
   949 => (x"71",x"87",x"f1",x"05"),
   950 => (x"0e",x"4f",x"26",x"48"),
   951 => (x"0e",x"5c",x"5b",x"5e"),
   952 => (x"4c",x"c0",x"4b",x"71"),
   953 => (x"70",x"87",x"f0",x"fe"),
   954 => (x"c0",x"02",x"99",x"49"),
   955 => (x"ec",x"c0",x"87",x"f9"),
   956 => (x"f2",x"c0",x"02",x"a9"),
   957 => (x"a9",x"fb",x"c0",x"87"),
   958 => (x"87",x"eb",x"c0",x"02"),
   959 => (x"ac",x"b7",x"66",x"cc"),
   960 => (x"d0",x"87",x"c7",x"03"),
   961 => (x"87",x"c2",x"02",x"66"),
   962 => (x"99",x"71",x"53",x"71"),
   963 => (x"c1",x"87",x"c2",x"02"),
   964 => (x"87",x"c3",x"fe",x"84"),
   965 => (x"02",x"99",x"49",x"70"),
   966 => (x"ec",x"c0",x"87",x"cd"),
   967 => (x"87",x"c7",x"02",x"a9"),
   968 => (x"05",x"a9",x"fb",x"c0"),
   969 => (x"d0",x"87",x"d5",x"ff"),
   970 => (x"87",x"c3",x"02",x"66"),
   971 => (x"c0",x"7b",x"97",x"c0"),
   972 => (x"c4",x"05",x"a9",x"ec"),
   973 => (x"c5",x"4a",x"74",x"87"),
   974 => (x"c0",x"4a",x"74",x"87"),
   975 => (x"48",x"72",x"8a",x"0a"),
   976 => (x"4d",x"26",x"87",x"c2"),
   977 => (x"4b",x"26",x"4c",x"26"),
   978 => (x"fd",x"1e",x"4f",x"26"),
   979 => (x"49",x"70",x"87",x"c9"),
   980 => (x"a9",x"b7",x"f0",x"c0"),
   981 => (x"c0",x"87",x"ca",x"04"),
   982 => (x"01",x"a9",x"b7",x"f9"),
   983 => (x"f0",x"c0",x"87",x"c3"),
   984 => (x"b7",x"c1",x"c1",x"89"),
   985 => (x"87",x"ca",x"04",x"a9"),
   986 => (x"a9",x"b7",x"da",x"c1"),
   987 => (x"c0",x"87",x"c3",x"01"),
   988 => (x"48",x"71",x"89",x"f7"),
   989 => (x"5e",x"0e",x"4f",x"26"),
   990 => (x"71",x"0e",x"5c",x"5b"),
   991 => (x"4c",x"d4",x"ff",x"4a"),
   992 => (x"ea",x"c0",x"49",x"72"),
   993 => (x"9b",x"4b",x"70",x"87"),
   994 => (x"c1",x"87",x"c2",x"02"),
   995 => (x"48",x"d0",x"ff",x"8b"),
   996 => (x"c1",x"78",x"c5",x"c8"),
   997 => (x"49",x"73",x"7c",x"d5"),
   998 => (x"e2",x"c2",x"31",x"c6"),
   999 => (x"4a",x"bf",x"97",x"df"),
  1000 => (x"70",x"b0",x"71",x"48"),
  1001 => (x"48",x"d0",x"ff",x"7c"),
  1002 => (x"48",x"73",x"78",x"c4"),
  1003 => (x"0e",x"87",x"d5",x"fe"),
  1004 => (x"5d",x"5c",x"5b",x"5e"),
  1005 => (x"71",x"86",x"f8",x"0e"),
  1006 => (x"fb",x"7e",x"c0",x"4c"),
  1007 => (x"4b",x"c0",x"87",x"e4"),
  1008 => (x"97",x"dc",x"c1",x"c1"),
  1009 => (x"a9",x"c0",x"49",x"bf"),
  1010 => (x"fb",x"87",x"cf",x"04"),
  1011 => (x"83",x"c1",x"87",x"f9"),
  1012 => (x"97",x"dc",x"c1",x"c1"),
  1013 => (x"06",x"ab",x"49",x"bf"),
  1014 => (x"c1",x"c1",x"87",x"f1"),
  1015 => (x"02",x"bf",x"97",x"dc"),
  1016 => (x"f2",x"fa",x"87",x"cf"),
  1017 => (x"99",x"49",x"70",x"87"),
  1018 => (x"c0",x"87",x"c6",x"02"),
  1019 => (x"f1",x"05",x"a9",x"ec"),
  1020 => (x"fa",x"4b",x"c0",x"87"),
  1021 => (x"4d",x"70",x"87",x"e1"),
  1022 => (x"c8",x"87",x"dc",x"fa"),
  1023 => (x"d6",x"fa",x"58",x"a6"),
  1024 => (x"c1",x"4a",x"70",x"87"),
  1025 => (x"49",x"a4",x"c8",x"83"),
  1026 => (x"ad",x"49",x"69",x"97"),
  1027 => (x"c0",x"87",x"c7",x"02"),
  1028 => (x"c0",x"05",x"ad",x"ff"),
  1029 => (x"a4",x"c9",x"87",x"e7"),
  1030 => (x"49",x"69",x"97",x"49"),
  1031 => (x"02",x"a9",x"66",x"c4"),
  1032 => (x"c0",x"48",x"87",x"c7"),
  1033 => (x"d4",x"05",x"a8",x"ff"),
  1034 => (x"49",x"a4",x"ca",x"87"),
  1035 => (x"aa",x"49",x"69",x"97"),
  1036 => (x"c0",x"87",x"c6",x"02"),
  1037 => (x"c4",x"05",x"aa",x"ff"),
  1038 => (x"d0",x"7e",x"c1",x"87"),
  1039 => (x"ad",x"ec",x"c0",x"87"),
  1040 => (x"c0",x"87",x"c6",x"02"),
  1041 => (x"c4",x"05",x"ad",x"fb"),
  1042 => (x"c1",x"4b",x"c0",x"87"),
  1043 => (x"fe",x"02",x"6e",x"7e"),
  1044 => (x"e9",x"f9",x"87",x"e1"),
  1045 => (x"f8",x"48",x"73",x"87"),
  1046 => (x"87",x"e6",x"fb",x"8e"),
  1047 => (x"5b",x"5e",x"0e",x"00"),
  1048 => (x"1e",x"0e",x"5d",x"5c"),
  1049 => (x"4c",x"c0",x"4b",x"71"),
  1050 => (x"c0",x"04",x"ab",x"4d"),
  1051 => (x"fe",x"c0",x"87",x"e8"),
  1052 => (x"9d",x"75",x"1e",x"ef"),
  1053 => (x"c0",x"87",x"c4",x"02"),
  1054 => (x"c1",x"87",x"c2",x"4a"),
  1055 => (x"f0",x"49",x"72",x"4a"),
  1056 => (x"86",x"c4",x"87",x"df"),
  1057 => (x"84",x"c1",x"7e",x"70"),
  1058 => (x"87",x"c2",x"05",x"6e"),
  1059 => (x"85",x"c1",x"4c",x"73"),
  1060 => (x"ff",x"06",x"ac",x"73"),
  1061 => (x"48",x"6e",x"87",x"d8"),
  1062 => (x"26",x"4d",x"26",x"26"),
  1063 => (x"26",x"4b",x"26",x"4c"),
  1064 => (x"5b",x"5e",x"0e",x"4f"),
  1065 => (x"1e",x"0e",x"5d",x"5c"),
  1066 => (x"de",x"49",x"4c",x"71"),
  1067 => (x"c1",x"f1",x"c2",x"91"),
  1068 => (x"97",x"85",x"71",x"4d"),
  1069 => (x"dd",x"c1",x"02",x"6d"),
  1070 => (x"ec",x"f0",x"c2",x"87"),
  1071 => (x"82",x"74",x"4a",x"bf"),
  1072 => (x"d8",x"fe",x"49",x"72"),
  1073 => (x"6e",x"7e",x"70",x"87"),
  1074 => (x"87",x"f3",x"c0",x"02"),
  1075 => (x"4b",x"f4",x"f0",x"c2"),
  1076 => (x"49",x"cb",x"4a",x"6e"),
  1077 => (x"87",x"d0",x"ff",x"fe"),
  1078 => (x"93",x"cb",x"4b",x"74"),
  1079 => (x"83",x"ca",x"e5",x"c1"),
  1080 => (x"c4",x"c1",x"83",x"c4"),
  1081 => (x"49",x"74",x"7b",x"da"),
  1082 => (x"87",x"c5",x"c3",x"c1"),
  1083 => (x"f1",x"c2",x"7b",x"75"),
  1084 => (x"49",x"bf",x"97",x"c0"),
  1085 => (x"f4",x"f0",x"c2",x"1e"),
  1086 => (x"e4",x"dd",x"c1",x"49"),
  1087 => (x"74",x"86",x"c4",x"87"),
  1088 => (x"ec",x"c2",x"c1",x"49"),
  1089 => (x"c1",x"49",x"c0",x"87"),
  1090 => (x"c2",x"87",x"cb",x"c4"),
  1091 => (x"c0",x"48",x"e8",x"f0"),
  1092 => (x"dd",x"49",x"c1",x"78"),
  1093 => (x"fd",x"26",x"87",x"cb"),
  1094 => (x"6f",x"4c",x"87",x"ff"),
  1095 => (x"6e",x"69",x"64",x"61"),
  1096 => (x"2e",x"2e",x"2e",x"67"),
  1097 => (x"5b",x"5e",x"0e",x"00"),
  1098 => (x"4b",x"71",x"0e",x"5c"),
  1099 => (x"ec",x"f0",x"c2",x"4a"),
  1100 => (x"49",x"72",x"82",x"bf"),
  1101 => (x"70",x"87",x"e6",x"fc"),
  1102 => (x"c4",x"02",x"9c",x"4c"),
  1103 => (x"e8",x"ec",x"49",x"87"),
  1104 => (x"ec",x"f0",x"c2",x"87"),
  1105 => (x"c1",x"78",x"c0",x"48"),
  1106 => (x"87",x"d5",x"dc",x"49"),
  1107 => (x"0e",x"87",x"cc",x"fd"),
  1108 => (x"5d",x"5c",x"5b",x"5e"),
  1109 => (x"c2",x"86",x"f4",x"0e"),
  1110 => (x"c0",x"4d",x"f6",x"e3"),
  1111 => (x"48",x"a6",x"c4",x"4c"),
  1112 => (x"f0",x"c2",x"78",x"c0"),
  1113 => (x"c0",x"49",x"bf",x"ec"),
  1114 => (x"c1",x"c1",x"06",x"a9"),
  1115 => (x"f6",x"e3",x"c2",x"87"),
  1116 => (x"c0",x"02",x"98",x"48"),
  1117 => (x"fe",x"c0",x"87",x"f8"),
  1118 => (x"66",x"c8",x"1e",x"ef"),
  1119 => (x"c4",x"87",x"c7",x"02"),
  1120 => (x"78",x"c0",x"48",x"a6"),
  1121 => (x"a6",x"c4",x"87",x"c5"),
  1122 => (x"c4",x"78",x"c1",x"48"),
  1123 => (x"d0",x"ec",x"49",x"66"),
  1124 => (x"70",x"86",x"c4",x"87"),
  1125 => (x"c4",x"84",x"c1",x"4d"),
  1126 => (x"80",x"c1",x"48",x"66"),
  1127 => (x"c2",x"58",x"a6",x"c8"),
  1128 => (x"49",x"bf",x"ec",x"f0"),
  1129 => (x"87",x"c6",x"03",x"ac"),
  1130 => (x"ff",x"05",x"9d",x"75"),
  1131 => (x"4c",x"c0",x"87",x"c8"),
  1132 => (x"c3",x"02",x"9d",x"75"),
  1133 => (x"fe",x"c0",x"87",x"e0"),
  1134 => (x"66",x"c8",x"1e",x"ef"),
  1135 => (x"cc",x"87",x"c7",x"02"),
  1136 => (x"78",x"c0",x"48",x"a6"),
  1137 => (x"a6",x"cc",x"87",x"c5"),
  1138 => (x"cc",x"78",x"c1",x"48"),
  1139 => (x"d0",x"eb",x"49",x"66"),
  1140 => (x"70",x"86",x"c4",x"87"),
  1141 => (x"c2",x"02",x"6e",x"7e"),
  1142 => (x"49",x"6e",x"87",x"e9"),
  1143 => (x"69",x"97",x"81",x"cb"),
  1144 => (x"02",x"99",x"d0",x"49"),
  1145 => (x"c1",x"87",x"d6",x"c1"),
  1146 => (x"74",x"4a",x"e5",x"c4"),
  1147 => (x"c1",x"91",x"cb",x"49"),
  1148 => (x"72",x"81",x"ca",x"e5"),
  1149 => (x"c3",x"81",x"c8",x"79"),
  1150 => (x"49",x"74",x"51",x"ff"),
  1151 => (x"f1",x"c2",x"91",x"de"),
  1152 => (x"85",x"71",x"4d",x"c1"),
  1153 => (x"7d",x"97",x"c1",x"c2"),
  1154 => (x"c0",x"49",x"a5",x"c1"),
  1155 => (x"ec",x"c2",x"51",x"e0"),
  1156 => (x"02",x"bf",x"97",x"c6"),
  1157 => (x"84",x"c1",x"87",x"d2"),
  1158 => (x"c2",x"4b",x"a5",x"c2"),
  1159 => (x"db",x"4a",x"c6",x"ec"),
  1160 => (x"c3",x"fa",x"fe",x"49"),
  1161 => (x"87",x"db",x"c1",x"87"),
  1162 => (x"c0",x"49",x"a5",x"cd"),
  1163 => (x"c2",x"84",x"c1",x"51"),
  1164 => (x"4a",x"6e",x"4b",x"a5"),
  1165 => (x"f9",x"fe",x"49",x"cb"),
  1166 => (x"c6",x"c1",x"87",x"ee"),
  1167 => (x"e1",x"c2",x"c1",x"87"),
  1168 => (x"cb",x"49",x"74",x"4a"),
  1169 => (x"ca",x"e5",x"c1",x"91"),
  1170 => (x"c2",x"79",x"72",x"81"),
  1171 => (x"bf",x"97",x"c6",x"ec"),
  1172 => (x"74",x"87",x"d8",x"02"),
  1173 => (x"c1",x"91",x"de",x"49"),
  1174 => (x"c1",x"f1",x"c2",x"84"),
  1175 => (x"c2",x"83",x"71",x"4b"),
  1176 => (x"dd",x"4a",x"c6",x"ec"),
  1177 => (x"ff",x"f8",x"fe",x"49"),
  1178 => (x"74",x"87",x"d8",x"87"),
  1179 => (x"c2",x"93",x"de",x"4b"),
  1180 => (x"cb",x"83",x"c1",x"f1"),
  1181 => (x"51",x"c0",x"49",x"a3"),
  1182 => (x"6e",x"73",x"84",x"c1"),
  1183 => (x"fe",x"49",x"cb",x"4a"),
  1184 => (x"c4",x"87",x"e5",x"f8"),
  1185 => (x"80",x"c1",x"48",x"66"),
  1186 => (x"c7",x"58",x"a6",x"c8"),
  1187 => (x"c5",x"c0",x"03",x"ac"),
  1188 => (x"fc",x"05",x"6e",x"87"),
  1189 => (x"48",x"74",x"87",x"e0"),
  1190 => (x"fc",x"f7",x"8e",x"f4"),
  1191 => (x"1e",x"73",x"1e",x"87"),
  1192 => (x"cb",x"49",x"4b",x"71"),
  1193 => (x"ca",x"e5",x"c1",x"91"),
  1194 => (x"4a",x"a1",x"c8",x"81"),
  1195 => (x"48",x"df",x"e2",x"c2"),
  1196 => (x"a1",x"c9",x"50",x"12"),
  1197 => (x"dc",x"c1",x"c1",x"4a"),
  1198 => (x"ca",x"50",x"12",x"48"),
  1199 => (x"c0",x"f1",x"c2",x"81"),
  1200 => (x"c2",x"50",x"11",x"48"),
  1201 => (x"bf",x"97",x"c0",x"f1"),
  1202 => (x"49",x"c0",x"1e",x"49"),
  1203 => (x"87",x"d1",x"d6",x"c1"),
  1204 => (x"48",x"e8",x"f0",x"c2"),
  1205 => (x"49",x"c1",x"78",x"de"),
  1206 => (x"26",x"87",x"c6",x"d6"),
  1207 => (x"1e",x"87",x"fe",x"f6"),
  1208 => (x"cb",x"49",x"4a",x"71"),
  1209 => (x"ca",x"e5",x"c1",x"91"),
  1210 => (x"11",x"81",x"c8",x"81"),
  1211 => (x"ec",x"f0",x"c2",x"48"),
  1212 => (x"ec",x"f0",x"c2",x"58"),
  1213 => (x"c1",x"78",x"c0",x"48"),
  1214 => (x"87",x"e5",x"d5",x"49"),
  1215 => (x"c0",x"1e",x"4f",x"26"),
  1216 => (x"d1",x"fc",x"c0",x"49"),
  1217 => (x"1e",x"4f",x"26",x"87"),
  1218 => (x"d2",x"02",x"99",x"71"),
  1219 => (x"df",x"e6",x"c1",x"87"),
  1220 => (x"f7",x"50",x"c0",x"48"),
  1221 => (x"df",x"cb",x"c1",x"80"),
  1222 => (x"c3",x"e5",x"c1",x"40"),
  1223 => (x"c1",x"87",x"ce",x"78"),
  1224 => (x"c1",x"48",x"db",x"e6"),
  1225 => (x"fc",x"78",x"fc",x"e4"),
  1226 => (x"fe",x"cb",x"c1",x"80"),
  1227 => (x"0e",x"4f",x"26",x"78"),
  1228 => (x"0e",x"5c",x"5b",x"5e"),
  1229 => (x"cb",x"4a",x"4c",x"71"),
  1230 => (x"ca",x"e5",x"c1",x"92"),
  1231 => (x"49",x"a2",x"c8",x"82"),
  1232 => (x"97",x"4b",x"a2",x"c9"),
  1233 => (x"97",x"1e",x"4b",x"6b"),
  1234 => (x"ca",x"1e",x"49",x"69"),
  1235 => (x"c0",x"49",x"12",x"82"),
  1236 => (x"c0",x"87",x"cc",x"e7"),
  1237 => (x"87",x"c9",x"d4",x"49"),
  1238 => (x"f9",x"c0",x"49",x"74"),
  1239 => (x"8e",x"f8",x"87",x"d3"),
  1240 => (x"1e",x"87",x"f8",x"f4"),
  1241 => (x"4b",x"71",x"1e",x"73"),
  1242 => (x"87",x"c3",x"ff",x"49"),
  1243 => (x"fe",x"fe",x"49",x"73"),
  1244 => (x"87",x"e9",x"f4",x"87"),
  1245 => (x"71",x"1e",x"73",x"1e"),
  1246 => (x"4a",x"a3",x"c6",x"4b"),
  1247 => (x"c1",x"87",x"db",x"02"),
  1248 => (x"87",x"d6",x"02",x"8a"),
  1249 => (x"da",x"c1",x"02",x"8a"),
  1250 => (x"c0",x"02",x"8a",x"87"),
  1251 => (x"02",x"8a",x"87",x"fc"),
  1252 => (x"8a",x"87",x"e1",x"c0"),
  1253 => (x"c1",x"87",x"cb",x"02"),
  1254 => (x"49",x"c7",x"87",x"db"),
  1255 => (x"c1",x"87",x"c0",x"fd"),
  1256 => (x"f0",x"c2",x"87",x"de"),
  1257 => (x"c1",x"02",x"bf",x"ec"),
  1258 => (x"c1",x"48",x"87",x"cb"),
  1259 => (x"f0",x"f0",x"c2",x"88"),
  1260 => (x"87",x"c1",x"c1",x"58"),
  1261 => (x"bf",x"f0",x"f0",x"c2"),
  1262 => (x"87",x"f9",x"c0",x"02"),
  1263 => (x"bf",x"ec",x"f0",x"c2"),
  1264 => (x"c2",x"80",x"c1",x"48"),
  1265 => (x"c0",x"58",x"f0",x"f0"),
  1266 => (x"f0",x"c2",x"87",x"eb"),
  1267 => (x"c6",x"49",x"bf",x"ec"),
  1268 => (x"f0",x"f0",x"c2",x"89"),
  1269 => (x"a9",x"b7",x"c0",x"59"),
  1270 => (x"c2",x"87",x"da",x"03"),
  1271 => (x"c0",x"48",x"ec",x"f0"),
  1272 => (x"c2",x"87",x"d2",x"78"),
  1273 => (x"02",x"bf",x"f0",x"f0"),
  1274 => (x"f0",x"c2",x"87",x"cb"),
  1275 => (x"c6",x"48",x"bf",x"ec"),
  1276 => (x"f0",x"f0",x"c2",x"80"),
  1277 => (x"d1",x"49",x"c0",x"58"),
  1278 => (x"49",x"73",x"87",x"e7"),
  1279 => (x"87",x"f1",x"f6",x"c0"),
  1280 => (x"0e",x"87",x"da",x"f2"),
  1281 => (x"0e",x"5c",x"5b",x"5e"),
  1282 => (x"66",x"cc",x"4c",x"71"),
  1283 => (x"cb",x"4b",x"74",x"1e"),
  1284 => (x"ca",x"e5",x"c1",x"93"),
  1285 => (x"4a",x"a3",x"c4",x"83"),
  1286 => (x"f2",x"fe",x"49",x"6a"),
  1287 => (x"ca",x"c1",x"87",x"da"),
  1288 => (x"a3",x"c8",x"7b",x"dd"),
  1289 => (x"51",x"66",x"d4",x"49"),
  1290 => (x"d8",x"49",x"a3",x"c9"),
  1291 => (x"a3",x"ca",x"51",x"66"),
  1292 => (x"51",x"66",x"dc",x"49"),
  1293 => (x"87",x"e3",x"f1",x"26"),
  1294 => (x"5c",x"5b",x"5e",x"0e"),
  1295 => (x"d0",x"ff",x"0e",x"5d"),
  1296 => (x"59",x"a6",x"d8",x"86"),
  1297 => (x"c0",x"48",x"a6",x"c4"),
  1298 => (x"c1",x"80",x"c4",x"78"),
  1299 => (x"c4",x"78",x"66",x"c4"),
  1300 => (x"c4",x"78",x"c1",x"80"),
  1301 => (x"c2",x"78",x"c1",x"80"),
  1302 => (x"c1",x"48",x"f0",x"f0"),
  1303 => (x"e8",x"f0",x"c2",x"78"),
  1304 => (x"a8",x"de",x"48",x"bf"),
  1305 => (x"f3",x"87",x"cb",x"05"),
  1306 => (x"49",x"70",x"87",x"e5"),
  1307 => (x"ce",x"59",x"a6",x"c8"),
  1308 => (x"ed",x"e8",x"87",x"f8"),
  1309 => (x"87",x"cf",x"e9",x"87"),
  1310 => (x"70",x"87",x"dc",x"e8"),
  1311 => (x"ac",x"fb",x"c0",x"4c"),
  1312 => (x"87",x"d0",x"c1",x"02"),
  1313 => (x"c1",x"05",x"66",x"d4"),
  1314 => (x"1e",x"c0",x"87",x"c2"),
  1315 => (x"c1",x"1e",x"c1",x"1e"),
  1316 => (x"c0",x"1e",x"fd",x"e6"),
  1317 => (x"87",x"eb",x"fd",x"49"),
  1318 => (x"4a",x"66",x"d0",x"c1"),
  1319 => (x"49",x"6a",x"82",x"c4"),
  1320 => (x"51",x"74",x"81",x"c7"),
  1321 => (x"1e",x"d8",x"1e",x"c1"),
  1322 => (x"81",x"c8",x"49",x"6a"),
  1323 => (x"d8",x"87",x"ec",x"e8"),
  1324 => (x"66",x"c4",x"c1",x"86"),
  1325 => (x"01",x"a8",x"c0",x"48"),
  1326 => (x"a6",x"c4",x"87",x"c7"),
  1327 => (x"ce",x"78",x"c1",x"48"),
  1328 => (x"66",x"c4",x"c1",x"87"),
  1329 => (x"cc",x"88",x"c1",x"48"),
  1330 => (x"87",x"c3",x"58",x"a6"),
  1331 => (x"cc",x"87",x"f8",x"e7"),
  1332 => (x"78",x"c2",x"48",x"a6"),
  1333 => (x"cd",x"02",x"9c",x"74"),
  1334 => (x"66",x"c4",x"87",x"cc"),
  1335 => (x"66",x"c8",x"c1",x"48"),
  1336 => (x"c1",x"cd",x"03",x"a8"),
  1337 => (x"48",x"a6",x"d8",x"87"),
  1338 => (x"ea",x"e6",x"78",x"c0"),
  1339 => (x"c1",x"4c",x"70",x"87"),
  1340 => (x"c2",x"05",x"ac",x"d0"),
  1341 => (x"66",x"d8",x"87",x"d6"),
  1342 => (x"87",x"ce",x"e9",x"7e"),
  1343 => (x"a6",x"dc",x"49",x"70"),
  1344 => (x"87",x"d3",x"e6",x"59"),
  1345 => (x"ec",x"c0",x"4c",x"70"),
  1346 => (x"ea",x"c1",x"05",x"ac"),
  1347 => (x"49",x"66",x"c4",x"87"),
  1348 => (x"c0",x"c1",x"91",x"cb"),
  1349 => (x"a1",x"c4",x"81",x"66"),
  1350 => (x"c8",x"4d",x"6a",x"4a"),
  1351 => (x"66",x"d8",x"4a",x"a1"),
  1352 => (x"df",x"cb",x"c1",x"52"),
  1353 => (x"87",x"ef",x"e5",x"79"),
  1354 => (x"02",x"9c",x"4c",x"70"),
  1355 => (x"fb",x"c0",x"87",x"d8"),
  1356 => (x"87",x"d2",x"02",x"ac"),
  1357 => (x"de",x"e5",x"55",x"74"),
  1358 => (x"9c",x"4c",x"70",x"87"),
  1359 => (x"c0",x"87",x"c7",x"02"),
  1360 => (x"ff",x"05",x"ac",x"fb"),
  1361 => (x"e0",x"c0",x"87",x"ee"),
  1362 => (x"55",x"c1",x"c2",x"55"),
  1363 => (x"d4",x"7d",x"97",x"c0"),
  1364 => (x"a9",x"6e",x"49",x"66"),
  1365 => (x"c4",x"87",x"db",x"05"),
  1366 => (x"66",x"c8",x"48",x"66"),
  1367 => (x"87",x"ca",x"04",x"a8"),
  1368 => (x"c1",x"48",x"66",x"c4"),
  1369 => (x"58",x"a6",x"c8",x"80"),
  1370 => (x"66",x"c8",x"87",x"c8"),
  1371 => (x"cc",x"88",x"c1",x"48"),
  1372 => (x"e2",x"e4",x"58",x"a6"),
  1373 => (x"c1",x"4c",x"70",x"87"),
  1374 => (x"c8",x"05",x"ac",x"d0"),
  1375 => (x"48",x"66",x"d0",x"87"),
  1376 => (x"a6",x"d4",x"80",x"c1"),
  1377 => (x"ac",x"d0",x"c1",x"58"),
  1378 => (x"87",x"ea",x"fd",x"02"),
  1379 => (x"d4",x"48",x"a6",x"dc"),
  1380 => (x"66",x"d8",x"78",x"66"),
  1381 => (x"a8",x"66",x"dc",x"48"),
  1382 => (x"87",x"dc",x"c9",x"05"),
  1383 => (x"48",x"a6",x"e0",x"c0"),
  1384 => (x"c4",x"78",x"f0",x"c0"),
  1385 => (x"78",x"66",x"cc",x"80"),
  1386 => (x"78",x"c0",x"80",x"c4"),
  1387 => (x"c0",x"48",x"74",x"7e"),
  1388 => (x"f0",x"c0",x"88",x"fb"),
  1389 => (x"98",x"70",x"58",x"a6"),
  1390 => (x"87",x"d7",x"c8",x"02"),
  1391 => (x"c0",x"88",x"cb",x"48"),
  1392 => (x"70",x"58",x"a6",x"f0"),
  1393 => (x"e9",x"c0",x"02",x"98"),
  1394 => (x"88",x"c9",x"48",x"87"),
  1395 => (x"58",x"a6",x"f0",x"c0"),
  1396 => (x"c3",x"02",x"98",x"70"),
  1397 => (x"c4",x"48",x"87",x"e1"),
  1398 => (x"a6",x"f0",x"c0",x"88"),
  1399 => (x"02",x"98",x"70",x"58"),
  1400 => (x"c1",x"48",x"87",x"de"),
  1401 => (x"a6",x"f0",x"c0",x"88"),
  1402 => (x"02",x"98",x"70",x"58"),
  1403 => (x"c7",x"87",x"c8",x"c3"),
  1404 => (x"e0",x"c0",x"87",x"db"),
  1405 => (x"78",x"c0",x"48",x"a6"),
  1406 => (x"c1",x"48",x"66",x"cc"),
  1407 => (x"58",x"a6",x"d0",x"80"),
  1408 => (x"70",x"87",x"d4",x"e2"),
  1409 => (x"ac",x"ec",x"c0",x"4c"),
  1410 => (x"c0",x"87",x"d5",x"02"),
  1411 => (x"c6",x"02",x"66",x"e0"),
  1412 => (x"a6",x"e4",x"c0",x"87"),
  1413 => (x"74",x"87",x"c9",x"5c"),
  1414 => (x"88",x"f0",x"c0",x"48"),
  1415 => (x"58",x"a6",x"e8",x"c0"),
  1416 => (x"02",x"ac",x"ec",x"c0"),
  1417 => (x"ee",x"e1",x"87",x"cc"),
  1418 => (x"c0",x"4c",x"70",x"87"),
  1419 => (x"ff",x"05",x"ac",x"ec"),
  1420 => (x"e0",x"c0",x"87",x"f4"),
  1421 => (x"66",x"d4",x"1e",x"66"),
  1422 => (x"ec",x"c0",x"1e",x"49"),
  1423 => (x"e6",x"c1",x"1e",x"66"),
  1424 => (x"66",x"d4",x"1e",x"fd"),
  1425 => (x"87",x"fb",x"f6",x"49"),
  1426 => (x"1e",x"ca",x"1e",x"c0"),
  1427 => (x"cb",x"49",x"66",x"dc"),
  1428 => (x"66",x"d8",x"c1",x"91"),
  1429 => (x"48",x"a6",x"d8",x"81"),
  1430 => (x"d8",x"78",x"a1",x"c4"),
  1431 => (x"e1",x"49",x"bf",x"66"),
  1432 => (x"86",x"d8",x"87",x"f9"),
  1433 => (x"06",x"a8",x"b7",x"c0"),
  1434 => (x"c1",x"87",x"c7",x"c1"),
  1435 => (x"c8",x"1e",x"de",x"1e"),
  1436 => (x"e1",x"49",x"bf",x"66"),
  1437 => (x"86",x"c8",x"87",x"e5"),
  1438 => (x"c0",x"48",x"49",x"70"),
  1439 => (x"e4",x"c0",x"88",x"08"),
  1440 => (x"b7",x"c0",x"58",x"a6"),
  1441 => (x"e9",x"c0",x"06",x"a8"),
  1442 => (x"66",x"e0",x"c0",x"87"),
  1443 => (x"a8",x"b7",x"dd",x"48"),
  1444 => (x"6e",x"87",x"df",x"03"),
  1445 => (x"e0",x"c0",x"49",x"bf"),
  1446 => (x"e0",x"c0",x"81",x"66"),
  1447 => (x"c1",x"49",x"66",x"51"),
  1448 => (x"81",x"bf",x"6e",x"81"),
  1449 => (x"c0",x"51",x"c1",x"c2"),
  1450 => (x"c2",x"49",x"66",x"e0"),
  1451 => (x"81",x"bf",x"6e",x"81"),
  1452 => (x"7e",x"c1",x"51",x"c0"),
  1453 => (x"e2",x"87",x"dc",x"c4"),
  1454 => (x"e4",x"c0",x"87",x"d0"),
  1455 => (x"c9",x"e2",x"58",x"a6"),
  1456 => (x"a6",x"e8",x"c0",x"87"),
  1457 => (x"a8",x"ec",x"c0",x"58"),
  1458 => (x"87",x"cb",x"c0",x"05"),
  1459 => (x"48",x"a6",x"e4",x"c0"),
  1460 => (x"78",x"66",x"e0",x"c0"),
  1461 => (x"ff",x"87",x"c4",x"c0"),
  1462 => (x"c4",x"87",x"fc",x"de"),
  1463 => (x"91",x"cb",x"49",x"66"),
  1464 => (x"48",x"66",x"c0",x"c1"),
  1465 => (x"7e",x"70",x"80",x"71"),
  1466 => (x"82",x"c8",x"4a",x"6e"),
  1467 => (x"81",x"ca",x"49",x"6e"),
  1468 => (x"51",x"66",x"e0",x"c0"),
  1469 => (x"49",x"66",x"e4",x"c0"),
  1470 => (x"e0",x"c0",x"81",x"c1"),
  1471 => (x"48",x"c1",x"89",x"66"),
  1472 => (x"49",x"70",x"30",x"71"),
  1473 => (x"97",x"71",x"89",x"c1"),
  1474 => (x"dd",x"f4",x"c2",x"7a"),
  1475 => (x"e0",x"c0",x"49",x"bf"),
  1476 => (x"6a",x"97",x"29",x"66"),
  1477 => (x"98",x"71",x"48",x"4a"),
  1478 => (x"58",x"a6",x"f0",x"c0"),
  1479 => (x"81",x"c4",x"49",x"6e"),
  1480 => (x"66",x"dc",x"4d",x"69"),
  1481 => (x"a8",x"66",x"d8",x"48"),
  1482 => (x"87",x"c8",x"c0",x"02"),
  1483 => (x"c0",x"48",x"a6",x"d8"),
  1484 => (x"87",x"c5",x"c0",x"78"),
  1485 => (x"c1",x"48",x"a6",x"d8"),
  1486 => (x"1e",x"66",x"d8",x"78"),
  1487 => (x"75",x"1e",x"e0",x"c0"),
  1488 => (x"d6",x"de",x"ff",x"49"),
  1489 => (x"70",x"86",x"c8",x"87"),
  1490 => (x"ac",x"b7",x"c0",x"4c"),
  1491 => (x"87",x"d4",x"c1",x"06"),
  1492 => (x"e0",x"c0",x"85",x"74"),
  1493 => (x"75",x"89",x"74",x"49"),
  1494 => (x"de",x"e1",x"c1",x"4b"),
  1495 => (x"e5",x"fe",x"71",x"4a"),
  1496 => (x"85",x"c2",x"87",x"c6"),
  1497 => (x"48",x"66",x"e8",x"c0"),
  1498 => (x"ec",x"c0",x"80",x"c1"),
  1499 => (x"ec",x"c0",x"58",x"a6"),
  1500 => (x"81",x"c1",x"49",x"66"),
  1501 => (x"c0",x"02",x"a9",x"70"),
  1502 => (x"a6",x"d8",x"87",x"c8"),
  1503 => (x"c0",x"78",x"c0",x"48"),
  1504 => (x"a6",x"d8",x"87",x"c5"),
  1505 => (x"d8",x"78",x"c1",x"48"),
  1506 => (x"a4",x"c2",x"1e",x"66"),
  1507 => (x"48",x"e0",x"c0",x"49"),
  1508 => (x"49",x"70",x"88",x"71"),
  1509 => (x"ff",x"49",x"75",x"1e"),
  1510 => (x"c8",x"87",x"c0",x"dd"),
  1511 => (x"a8",x"b7",x"c0",x"86"),
  1512 => (x"87",x"c0",x"ff",x"01"),
  1513 => (x"02",x"66",x"e8",x"c0"),
  1514 => (x"6e",x"87",x"d1",x"c0"),
  1515 => (x"c0",x"81",x"c9",x"49"),
  1516 => (x"6e",x"51",x"66",x"e8"),
  1517 => (x"ef",x"cc",x"c1",x"48"),
  1518 => (x"87",x"cc",x"c0",x"78"),
  1519 => (x"81",x"c9",x"49",x"6e"),
  1520 => (x"48",x"6e",x"51",x"c2"),
  1521 => (x"78",x"e3",x"cd",x"c1"),
  1522 => (x"c6",x"c0",x"7e",x"c1"),
  1523 => (x"f6",x"db",x"ff",x"87"),
  1524 => (x"6e",x"4c",x"70",x"87"),
  1525 => (x"87",x"f5",x"c0",x"02"),
  1526 => (x"c8",x"48",x"66",x"c4"),
  1527 => (x"c0",x"04",x"a8",x"66"),
  1528 => (x"66",x"c4",x"87",x"cb"),
  1529 => (x"c8",x"80",x"c1",x"48"),
  1530 => (x"e0",x"c0",x"58",x"a6"),
  1531 => (x"48",x"66",x"c8",x"87"),
  1532 => (x"a6",x"cc",x"88",x"c1"),
  1533 => (x"87",x"d5",x"c0",x"58"),
  1534 => (x"05",x"ac",x"c6",x"c1"),
  1535 => (x"cc",x"87",x"c8",x"c0"),
  1536 => (x"80",x"c1",x"48",x"66"),
  1537 => (x"ff",x"58",x"a6",x"d0"),
  1538 => (x"70",x"87",x"fc",x"da"),
  1539 => (x"48",x"66",x"d0",x"4c"),
  1540 => (x"a6",x"d4",x"80",x"c1"),
  1541 => (x"02",x"9c",x"74",x"58"),
  1542 => (x"c4",x"87",x"cb",x"c0"),
  1543 => (x"c8",x"c1",x"48",x"66"),
  1544 => (x"f2",x"04",x"a8",x"66"),
  1545 => (x"da",x"ff",x"87",x"ff"),
  1546 => (x"66",x"c4",x"87",x"d4"),
  1547 => (x"03",x"a8",x"c7",x"48"),
  1548 => (x"c2",x"87",x"e5",x"c0"),
  1549 => (x"c0",x"48",x"f0",x"f0"),
  1550 => (x"49",x"66",x"c4",x"78"),
  1551 => (x"c0",x"c1",x"91",x"cb"),
  1552 => (x"a1",x"c4",x"81",x"66"),
  1553 => (x"c0",x"4a",x"6a",x"4a"),
  1554 => (x"66",x"c4",x"79",x"52"),
  1555 => (x"c8",x"80",x"c1",x"48"),
  1556 => (x"a8",x"c7",x"58",x"a6"),
  1557 => (x"87",x"db",x"ff",x"04"),
  1558 => (x"e0",x"8e",x"d0",x"ff"),
  1559 => (x"20",x"3a",x"87",x"fb"),
  1560 => (x"1e",x"73",x"1e",x"00"),
  1561 => (x"02",x"9b",x"4b",x"71"),
  1562 => (x"f0",x"c2",x"87",x"c6"),
  1563 => (x"78",x"c0",x"48",x"ec"),
  1564 => (x"f0",x"c2",x"1e",x"c7"),
  1565 => (x"1e",x"49",x"bf",x"ec"),
  1566 => (x"1e",x"ca",x"e5",x"c1"),
  1567 => (x"bf",x"e8",x"f0",x"c2"),
  1568 => (x"87",x"f4",x"ee",x"49"),
  1569 => (x"f0",x"c2",x"86",x"cc"),
  1570 => (x"e9",x"49",x"bf",x"e8"),
  1571 => (x"9b",x"73",x"87",x"f9"),
  1572 => (x"c1",x"87",x"c8",x"02"),
  1573 => (x"c0",x"49",x"ca",x"e5"),
  1574 => (x"ff",x"87",x"e8",x"e5"),
  1575 => (x"1e",x"87",x"fe",x"df"),
  1576 => (x"48",x"df",x"e2",x"c2"),
  1577 => (x"e6",x"c1",x"50",x"c0"),
  1578 => (x"c0",x"49",x"bf",x"ed"),
  1579 => (x"c0",x"87",x"c5",x"fb"),
  1580 => (x"1e",x"4f",x"26",x"48"),
  1581 => (x"c1",x"87",x"e5",x"c7"),
  1582 => (x"87",x"e5",x"fe",x"49"),
  1583 => (x"87",x"e0",x"e9",x"fe"),
  1584 => (x"cd",x"02",x"98",x"70"),
  1585 => (x"dd",x"f2",x"fe",x"87"),
  1586 => (x"02",x"98",x"70",x"87"),
  1587 => (x"4a",x"c1",x"87",x"c4"),
  1588 => (x"4a",x"c0",x"87",x"c2"),
  1589 => (x"ce",x"05",x"9a",x"72"),
  1590 => (x"c1",x"1e",x"c0",x"87"),
  1591 => (x"c0",x"49",x"c3",x"e4"),
  1592 => (x"c4",x"87",x"ef",x"f0"),
  1593 => (x"c0",x"87",x"fe",x"86"),
  1594 => (x"ce",x"e4",x"c1",x"1e"),
  1595 => (x"e1",x"f0",x"c0",x"49"),
  1596 => (x"fe",x"1e",x"c0",x"87"),
  1597 => (x"49",x"70",x"87",x"e9"),
  1598 => (x"87",x"d6",x"f0",x"c0"),
  1599 => (x"f8",x"87",x"dc",x"c3"),
  1600 => (x"53",x"4f",x"26",x"8e"),
  1601 => (x"61",x"66",x"20",x"44"),
  1602 => (x"64",x"65",x"6c",x"69"),
  1603 => (x"6f",x"42",x"00",x"2e"),
  1604 => (x"6e",x"69",x"74",x"6f"),
  1605 => (x"2e",x"2e",x"2e",x"67"),
  1606 => (x"e8",x"c0",x"1e",x"00"),
  1607 => (x"f3",x"c0",x"87",x"c1"),
  1608 => (x"87",x"f6",x"87",x"e6"),
  1609 => (x"c2",x"1e",x"4f",x"26"),
  1610 => (x"c0",x"48",x"ec",x"f0"),
  1611 => (x"e8",x"f0",x"c2",x"78"),
  1612 => (x"fd",x"78",x"c0",x"48"),
  1613 => (x"87",x"e1",x"87",x"fd"),
  1614 => (x"4f",x"26",x"48",x"c0"),
  1615 => (x"78",x"45",x"20",x"80"),
  1616 => (x"80",x"00",x"74",x"69"),
  1617 => (x"63",x"61",x"42",x"20"),
  1618 => (x"12",x"df",x"00",x"6b"),
  1619 => (x"2c",x"41",x"00",x"00"),
  1620 => (x"00",x"00",x"00",x"00"),
  1621 => (x"00",x"12",x"df",x"00"),
  1622 => (x"00",x"2c",x"5f",x"00"),
  1623 => (x"00",x"00",x"00",x"00"),
  1624 => (x"00",x"00",x"12",x"df"),
  1625 => (x"00",x"00",x"2c",x"7d"),
  1626 => (x"df",x"00",x"00",x"00"),
  1627 => (x"9b",x"00",x"00",x"12"),
  1628 => (x"00",x"00",x"00",x"2c"),
  1629 => (x"12",x"df",x"00",x"00"),
  1630 => (x"2c",x"b9",x"00",x"00"),
  1631 => (x"00",x"00",x"00",x"00"),
  1632 => (x"00",x"12",x"df",x"00"),
  1633 => (x"00",x"2c",x"d7",x"00"),
  1634 => (x"00",x"00",x"00",x"00"),
  1635 => (x"00",x"00",x"12",x"df"),
  1636 => (x"00",x"00",x"2c",x"f5"),
  1637 => (x"df",x"00",x"00",x"00"),
  1638 => (x"00",x"00",x"00",x"12"),
  1639 => (x"00",x"00",x"00",x"00"),
  1640 => (x"13",x"74",x"00",x"00"),
  1641 => (x"00",x"00",x"00",x"00"),
  1642 => (x"00",x"00",x"00",x"00"),
  1643 => (x"00",x"19",x"b1",x"00"),
  1644 => (x"4f",x"4f",x"42",x"00"),
  1645 => (x"20",x"20",x"20",x"54"),
  1646 => (x"4d",x"4f",x"52",x"20"),
  1647 => (x"61",x"6f",x"4c",x"00"),
  1648 => (x"2e",x"2a",x"20",x"64"),
  1649 => (x"f0",x"fe",x"1e",x"00"),
  1650 => (x"cd",x"78",x"c0",x"48"),
  1651 => (x"26",x"09",x"79",x"09"),
  1652 => (x"fe",x"1e",x"1e",x"4f"),
  1653 => (x"48",x"7e",x"bf",x"f0"),
  1654 => (x"1e",x"4f",x"26",x"26"),
  1655 => (x"c1",x"48",x"f0",x"fe"),
  1656 => (x"1e",x"4f",x"26",x"78"),
  1657 => (x"c0",x"48",x"f0",x"fe"),
  1658 => (x"1e",x"4f",x"26",x"78"),
  1659 => (x"52",x"c0",x"4a",x"71"),
  1660 => (x"0e",x"4f",x"26",x"52"),
  1661 => (x"5d",x"5c",x"5b",x"5e"),
  1662 => (x"71",x"86",x"f4",x"0e"),
  1663 => (x"7e",x"6d",x"97",x"4d"),
  1664 => (x"97",x"4c",x"a5",x"c1"),
  1665 => (x"a6",x"c8",x"48",x"6c"),
  1666 => (x"c4",x"48",x"6e",x"58"),
  1667 => (x"c5",x"05",x"a8",x"66"),
  1668 => (x"c0",x"48",x"ff",x"87"),
  1669 => (x"ca",x"ff",x"87",x"e6"),
  1670 => (x"49",x"a5",x"c2",x"87"),
  1671 => (x"71",x"4b",x"6c",x"97"),
  1672 => (x"6b",x"97",x"4b",x"a3"),
  1673 => (x"7e",x"6c",x"97",x"4b"),
  1674 => (x"80",x"c1",x"48",x"6e"),
  1675 => (x"c7",x"58",x"a6",x"c8"),
  1676 => (x"58",x"a6",x"cc",x"98"),
  1677 => (x"fe",x"7c",x"97",x"70"),
  1678 => (x"48",x"73",x"87",x"e1"),
  1679 => (x"4d",x"26",x"8e",x"f4"),
  1680 => (x"4b",x"26",x"4c",x"26"),
  1681 => (x"5e",x"0e",x"4f",x"26"),
  1682 => (x"f4",x"0e",x"5c",x"5b"),
  1683 => (x"d8",x"4c",x"71",x"86"),
  1684 => (x"ff",x"c3",x"4a",x"66"),
  1685 => (x"4b",x"a4",x"c2",x"9a"),
  1686 => (x"73",x"49",x"6c",x"97"),
  1687 => (x"51",x"72",x"49",x"a1"),
  1688 => (x"6e",x"7e",x"6c",x"97"),
  1689 => (x"c8",x"80",x"c1",x"48"),
  1690 => (x"98",x"c7",x"58",x"a6"),
  1691 => (x"70",x"58",x"a6",x"cc"),
  1692 => (x"ff",x"8e",x"f4",x"54"),
  1693 => (x"1e",x"1e",x"87",x"ca"),
  1694 => (x"e0",x"87",x"e8",x"fd"),
  1695 => (x"c0",x"49",x"4a",x"bf"),
  1696 => (x"02",x"99",x"c0",x"e0"),
  1697 => (x"1e",x"72",x"87",x"cb"),
  1698 => (x"49",x"d3",x"f4",x"c2"),
  1699 => (x"c4",x"87",x"f7",x"fe"),
  1700 => (x"87",x"fd",x"fc",x"86"),
  1701 => (x"c2",x"fd",x"7e",x"70"),
  1702 => (x"4f",x"26",x"26",x"87"),
  1703 => (x"d3",x"f4",x"c2",x"1e"),
  1704 => (x"87",x"c7",x"fd",x"49"),
  1705 => (x"49",x"f6",x"e9",x"c1"),
  1706 => (x"c5",x"87",x"da",x"fc"),
  1707 => (x"4f",x"26",x"87",x"d9"),
  1708 => (x"5c",x"5b",x"5e",x"0e"),
  1709 => (x"f4",x"c2",x"0e",x"5d"),
  1710 => (x"c1",x"4a",x"bf",x"f2"),
  1711 => (x"49",x"bf",x"c4",x"ec"),
  1712 => (x"71",x"bc",x"72",x"4c"),
  1713 => (x"87",x"db",x"fc",x"4d"),
  1714 => (x"49",x"74",x"4b",x"c0"),
  1715 => (x"d5",x"02",x"99",x"d0"),
  1716 => (x"d0",x"49",x"75",x"87"),
  1717 => (x"c0",x"1e",x"71",x"99"),
  1718 => (x"d6",x"f2",x"c1",x"1e"),
  1719 => (x"12",x"82",x"73",x"4a"),
  1720 => (x"87",x"e4",x"c0",x"49"),
  1721 => (x"2c",x"c1",x"86",x"c8"),
  1722 => (x"ab",x"c8",x"83",x"2d"),
  1723 => (x"87",x"da",x"ff",x"04"),
  1724 => (x"c1",x"87",x"e8",x"fb"),
  1725 => (x"c2",x"48",x"c4",x"ec"),
  1726 => (x"78",x"bf",x"f2",x"f4"),
  1727 => (x"4c",x"26",x"4d",x"26"),
  1728 => (x"4f",x"26",x"4b",x"26"),
  1729 => (x"00",x"00",x"00",x"00"),
  1730 => (x"48",x"d0",x"ff",x"1e"),
  1731 => (x"ff",x"78",x"e1",x"c8"),
  1732 => (x"78",x"c5",x"48",x"d4"),
  1733 => (x"c3",x"02",x"66",x"c4"),
  1734 => (x"78",x"e0",x"c3",x"87"),
  1735 => (x"c6",x"02",x"66",x"c8"),
  1736 => (x"48",x"d4",x"ff",x"87"),
  1737 => (x"ff",x"78",x"f0",x"c3"),
  1738 => (x"78",x"71",x"48",x"d4"),
  1739 => (x"c8",x"48",x"d0",x"ff"),
  1740 => (x"e0",x"c0",x"78",x"e1"),
  1741 => (x"0e",x"4f",x"26",x"78"),
  1742 => (x"0e",x"5c",x"5b",x"5e"),
  1743 => (x"f4",x"c2",x"4c",x"71"),
  1744 => (x"ee",x"fa",x"49",x"d3"),
  1745 => (x"c0",x"4a",x"70",x"87"),
  1746 => (x"c2",x"04",x"aa",x"b7"),
  1747 => (x"e0",x"c3",x"87",x"e3"),
  1748 => (x"87",x"c9",x"05",x"aa"),
  1749 => (x"48",x"fa",x"ef",x"c1"),
  1750 => (x"d4",x"c2",x"78",x"c1"),
  1751 => (x"aa",x"f0",x"c3",x"87"),
  1752 => (x"c1",x"87",x"c9",x"05"),
  1753 => (x"c1",x"48",x"f6",x"ef"),
  1754 => (x"87",x"f5",x"c1",x"78"),
  1755 => (x"bf",x"fa",x"ef",x"c1"),
  1756 => (x"72",x"87",x"c7",x"02"),
  1757 => (x"b3",x"c0",x"c2",x"4b"),
  1758 => (x"4b",x"72",x"87",x"c2"),
  1759 => (x"d1",x"05",x"9c",x"74"),
  1760 => (x"f6",x"ef",x"c1",x"87"),
  1761 => (x"ef",x"c1",x"1e",x"bf"),
  1762 => (x"72",x"1e",x"bf",x"fa"),
  1763 => (x"87",x"f8",x"fd",x"49"),
  1764 => (x"ef",x"c1",x"86",x"c8"),
  1765 => (x"c0",x"02",x"bf",x"f6"),
  1766 => (x"49",x"73",x"87",x"e0"),
  1767 => (x"91",x"29",x"b7",x"c4"),
  1768 => (x"81",x"d6",x"f1",x"c1"),
  1769 => (x"9a",x"cf",x"4a",x"73"),
  1770 => (x"48",x"c1",x"92",x"c2"),
  1771 => (x"4a",x"70",x"30",x"72"),
  1772 => (x"48",x"72",x"ba",x"ff"),
  1773 => (x"79",x"70",x"98",x"69"),
  1774 => (x"49",x"73",x"87",x"db"),
  1775 => (x"91",x"29",x"b7",x"c4"),
  1776 => (x"81",x"d6",x"f1",x"c1"),
  1777 => (x"9a",x"cf",x"4a",x"73"),
  1778 => (x"48",x"c3",x"92",x"c2"),
  1779 => (x"4a",x"70",x"30",x"72"),
  1780 => (x"70",x"b0",x"69",x"48"),
  1781 => (x"fa",x"ef",x"c1",x"79"),
  1782 => (x"c1",x"78",x"c0",x"48"),
  1783 => (x"c0",x"48",x"f6",x"ef"),
  1784 => (x"d3",x"f4",x"c2",x"78"),
  1785 => (x"87",x"cb",x"f8",x"49"),
  1786 => (x"b7",x"c0",x"4a",x"70"),
  1787 => (x"dd",x"fd",x"03",x"aa"),
  1788 => (x"fc",x"48",x"c0",x"87"),
  1789 => (x"00",x"00",x"87",x"c8"),
  1790 => (x"00",x"00",x"00",x"00"),
  1791 => (x"71",x"1e",x"00",x"00"),
  1792 => (x"f2",x"fc",x"49",x"4a"),
  1793 => (x"1e",x"4f",x"26",x"87"),
  1794 => (x"49",x"72",x"4a",x"c0"),
  1795 => (x"f1",x"c1",x"91",x"c4"),
  1796 => (x"79",x"c0",x"81",x"d6"),
  1797 => (x"b7",x"d0",x"82",x"c1"),
  1798 => (x"87",x"ee",x"04",x"aa"),
  1799 => (x"5e",x"0e",x"4f",x"26"),
  1800 => (x"0e",x"5d",x"5c",x"5b"),
  1801 => (x"fa",x"f6",x"4d",x"71"),
  1802 => (x"c4",x"4a",x"75",x"87"),
  1803 => (x"c1",x"92",x"2a",x"b7"),
  1804 => (x"75",x"82",x"d6",x"f1"),
  1805 => (x"c2",x"9c",x"cf",x"4c"),
  1806 => (x"4b",x"49",x"6a",x"94"),
  1807 => (x"9b",x"c3",x"2b",x"74"),
  1808 => (x"30",x"74",x"48",x"c2"),
  1809 => (x"bc",x"ff",x"4c",x"70"),
  1810 => (x"98",x"71",x"48",x"74"),
  1811 => (x"ca",x"f6",x"7a",x"70"),
  1812 => (x"fa",x"48",x"73",x"87"),
  1813 => (x"00",x"00",x"87",x"e6"),
  1814 => (x"00",x"00",x"00",x"00"),
  1815 => (x"00",x"00",x"00",x"00"),
  1816 => (x"00",x"00",x"00",x"00"),
  1817 => (x"00",x"00",x"00",x"00"),
  1818 => (x"00",x"00",x"00",x"00"),
  1819 => (x"00",x"00",x"00",x"00"),
  1820 => (x"00",x"00",x"00",x"00"),
  1821 => (x"00",x"00",x"00",x"00"),
  1822 => (x"00",x"00",x"00",x"00"),
  1823 => (x"00",x"00",x"00",x"00"),
  1824 => (x"00",x"00",x"00",x"00"),
  1825 => (x"00",x"00",x"00",x"00"),
  1826 => (x"00",x"00",x"00",x"00"),
  1827 => (x"00",x"00",x"00",x"00"),
  1828 => (x"00",x"00",x"00",x"00"),
  1829 => (x"1e",x"16",x"00",x"00"),
  1830 => (x"36",x"2e",x"25",x"26"),
  1831 => (x"ff",x"1e",x"3e",x"3d"),
  1832 => (x"e1",x"c8",x"48",x"d0"),
  1833 => (x"ff",x"48",x"71",x"78"),
  1834 => (x"26",x"78",x"08",x"d4"),
  1835 => (x"d0",x"ff",x"1e",x"4f"),
  1836 => (x"78",x"e1",x"c8",x"48"),
  1837 => (x"d4",x"ff",x"48",x"71"),
  1838 => (x"66",x"c4",x"78",x"08"),
  1839 => (x"08",x"d4",x"ff",x"48"),
  1840 => (x"1e",x"4f",x"26",x"78"),
  1841 => (x"66",x"c4",x"4a",x"71"),
  1842 => (x"49",x"72",x"1e",x"49"),
  1843 => (x"ff",x"87",x"de",x"ff"),
  1844 => (x"e0",x"c0",x"48",x"d0"),
  1845 => (x"4f",x"26",x"26",x"78"),
  1846 => (x"c2",x"4a",x"71",x"1e"),
  1847 => (x"c3",x"03",x"aa",x"b7"),
  1848 => (x"87",x"c2",x"82",x"87"),
  1849 => (x"66",x"c4",x"82",x"ce"),
  1850 => (x"ff",x"49",x"72",x"1e"),
  1851 => (x"26",x"26",x"87",x"d5"),
  1852 => (x"d4",x"ff",x"1e",x"4f"),
  1853 => (x"7a",x"ff",x"c3",x"4a"),
  1854 => (x"c8",x"48",x"d0",x"ff"),
  1855 => (x"7a",x"de",x"78",x"e1"),
  1856 => (x"bf",x"dd",x"f4",x"c2"),
  1857 => (x"c8",x"48",x"49",x"7a"),
  1858 => (x"71",x"7a",x"70",x"28"),
  1859 => (x"70",x"28",x"d0",x"48"),
  1860 => (x"d8",x"48",x"71",x"7a"),
  1861 => (x"ff",x"7a",x"70",x"28"),
  1862 => (x"e0",x"c0",x"48",x"d0"),
  1863 => (x"0e",x"4f",x"26",x"78"),
  1864 => (x"5d",x"5c",x"5b",x"5e"),
  1865 => (x"c2",x"4c",x"71",x"0e"),
  1866 => (x"4d",x"bf",x"dd",x"f4"),
  1867 => (x"d0",x"2b",x"74",x"4b"),
  1868 => (x"83",x"c1",x"9b",x"66"),
  1869 => (x"04",x"ab",x"66",x"d4"),
  1870 => (x"4b",x"c0",x"87",x"c2"),
  1871 => (x"66",x"d0",x"4a",x"74"),
  1872 => (x"ff",x"31",x"72",x"49"),
  1873 => (x"73",x"99",x"75",x"b9"),
  1874 => (x"70",x"30",x"72",x"48"),
  1875 => (x"b0",x"71",x"48",x"4a"),
  1876 => (x"58",x"e1",x"f4",x"c2"),
  1877 => (x"26",x"87",x"da",x"fe"),
  1878 => (x"26",x"4c",x"26",x"4d"),
  1879 => (x"1e",x"4f",x"26",x"4b"),
  1880 => (x"c8",x"48",x"d0",x"ff"),
  1881 => (x"48",x"71",x"78",x"c9"),
  1882 => (x"78",x"08",x"d4",x"ff"),
  1883 => (x"71",x"1e",x"4f",x"26"),
  1884 => (x"87",x"eb",x"49",x"4a"),
  1885 => (x"c8",x"48",x"d0",x"ff"),
  1886 => (x"1e",x"4f",x"26",x"78"),
  1887 => (x"4b",x"71",x"1e",x"73"),
  1888 => (x"bf",x"ed",x"f4",x"c2"),
  1889 => (x"c2",x"87",x"c3",x"02"),
  1890 => (x"d0",x"ff",x"87",x"eb"),
  1891 => (x"78",x"c9",x"c8",x"48"),
  1892 => (x"e0",x"c0",x"49",x"73"),
  1893 => (x"48",x"d4",x"ff",x"b1"),
  1894 => (x"f4",x"c2",x"78",x"71"),
  1895 => (x"78",x"c0",x"48",x"e1"),
  1896 => (x"c5",x"02",x"66",x"c8"),
  1897 => (x"49",x"ff",x"c3",x"87"),
  1898 => (x"49",x"c0",x"87",x"c2"),
  1899 => (x"59",x"e9",x"f4",x"c2"),
  1900 => (x"c6",x"02",x"66",x"cc"),
  1901 => (x"d5",x"d5",x"c5",x"87"),
  1902 => (x"cf",x"87",x"c4",x"4a"),
  1903 => (x"c2",x"4a",x"ff",x"ff"),
  1904 => (x"c2",x"5a",x"ed",x"f4"),
  1905 => (x"c1",x"48",x"ed",x"f4"),
  1906 => (x"26",x"87",x"c4",x"78"),
  1907 => (x"26",x"4c",x"26",x"4d"),
  1908 => (x"0e",x"4f",x"26",x"4b"),
  1909 => (x"5d",x"5c",x"5b",x"5e"),
  1910 => (x"c2",x"4a",x"71",x"0e"),
  1911 => (x"4c",x"bf",x"e9",x"f4"),
  1912 => (x"cb",x"02",x"9a",x"72"),
  1913 => (x"91",x"c8",x"49",x"87"),
  1914 => (x"4b",x"f1",x"f5",x"c1"),
  1915 => (x"87",x"c4",x"83",x"71"),
  1916 => (x"4b",x"f1",x"f9",x"c1"),
  1917 => (x"49",x"13",x"4d",x"c0"),
  1918 => (x"f4",x"c2",x"99",x"74"),
  1919 => (x"ff",x"b9",x"bf",x"e5"),
  1920 => (x"78",x"71",x"48",x"d4"),
  1921 => (x"85",x"2c",x"b7",x"c1"),
  1922 => (x"04",x"ad",x"b7",x"c8"),
  1923 => (x"f4",x"c2",x"87",x"e8"),
  1924 => (x"c8",x"48",x"bf",x"e1"),
  1925 => (x"e5",x"f4",x"c2",x"80"),
  1926 => (x"87",x"ef",x"fe",x"58"),
  1927 => (x"71",x"1e",x"73",x"1e"),
  1928 => (x"9a",x"4a",x"13",x"4b"),
  1929 => (x"72",x"87",x"cb",x"02"),
  1930 => (x"87",x"e7",x"fe",x"49"),
  1931 => (x"05",x"9a",x"4a",x"13"),
  1932 => (x"da",x"fe",x"87",x"f5"),
  1933 => (x"f4",x"c2",x"1e",x"87"),
  1934 => (x"c2",x"49",x"bf",x"e1"),
  1935 => (x"c1",x"48",x"e1",x"f4"),
  1936 => (x"c0",x"c4",x"78",x"a1"),
  1937 => (x"db",x"03",x"a9",x"b7"),
  1938 => (x"48",x"d4",x"ff",x"87"),
  1939 => (x"bf",x"e5",x"f4",x"c2"),
  1940 => (x"e1",x"f4",x"c2",x"78"),
  1941 => (x"f4",x"c2",x"49",x"bf"),
  1942 => (x"a1",x"c1",x"48",x"e1"),
  1943 => (x"b7",x"c0",x"c4",x"78"),
  1944 => (x"87",x"e5",x"04",x"a9"),
  1945 => (x"c8",x"48",x"d0",x"ff"),
  1946 => (x"ed",x"f4",x"c2",x"78"),
  1947 => (x"26",x"78",x"c0",x"48"),
  1948 => (x"00",x"00",x"00",x"4f"),
  1949 => (x"00",x"00",x"00",x"00"),
  1950 => (x"00",x"00",x"00",x"00"),
  1951 => (x"00",x"00",x"5f",x"5f"),
  1952 => (x"03",x"03",x"00",x"00"),
  1953 => (x"00",x"03",x"03",x"00"),
  1954 => (x"7f",x"7f",x"14",x"00"),
  1955 => (x"14",x"7f",x"7f",x"14"),
  1956 => (x"2e",x"24",x"00",x"00"),
  1957 => (x"12",x"3a",x"6b",x"6b"),
  1958 => (x"36",x"6a",x"4c",x"00"),
  1959 => (x"32",x"56",x"6c",x"18"),
  1960 => (x"4f",x"7e",x"30",x"00"),
  1961 => (x"68",x"3a",x"77",x"59"),
  1962 => (x"04",x"00",x"00",x"40"),
  1963 => (x"00",x"00",x"03",x"07"),
  1964 => (x"1c",x"00",x"00",x"00"),
  1965 => (x"00",x"41",x"63",x"3e"),
  1966 => (x"41",x"00",x"00",x"00"),
  1967 => (x"00",x"1c",x"3e",x"63"),
  1968 => (x"3e",x"2a",x"08",x"00"),
  1969 => (x"2a",x"3e",x"1c",x"1c"),
  1970 => (x"08",x"08",x"00",x"08"),
  1971 => (x"08",x"08",x"3e",x"3e"),
  1972 => (x"80",x"00",x"00",x"00"),
  1973 => (x"00",x"00",x"60",x"e0"),
  1974 => (x"08",x"08",x"00",x"00"),
  1975 => (x"08",x"08",x"08",x"08"),
  1976 => (x"00",x"00",x"00",x"00"),
  1977 => (x"00",x"00",x"60",x"60"),
  1978 => (x"30",x"60",x"40",x"00"),
  1979 => (x"03",x"06",x"0c",x"18"),
  1980 => (x"7f",x"3e",x"00",x"01"),
  1981 => (x"3e",x"7f",x"4d",x"59"),
  1982 => (x"06",x"04",x"00",x"00"),
  1983 => (x"00",x"00",x"7f",x"7f"),
  1984 => (x"63",x"42",x"00",x"00"),
  1985 => (x"46",x"4f",x"59",x"71"),
  1986 => (x"63",x"22",x"00",x"00"),
  1987 => (x"36",x"7f",x"49",x"49"),
  1988 => (x"16",x"1c",x"18",x"00"),
  1989 => (x"10",x"7f",x"7f",x"13"),
  1990 => (x"67",x"27",x"00",x"00"),
  1991 => (x"39",x"7d",x"45",x"45"),
  1992 => (x"7e",x"3c",x"00",x"00"),
  1993 => (x"30",x"79",x"49",x"4b"),
  1994 => (x"01",x"01",x"00",x"00"),
  1995 => (x"07",x"0f",x"79",x"71"),
  1996 => (x"7f",x"36",x"00",x"00"),
  1997 => (x"36",x"7f",x"49",x"49"),
  1998 => (x"4f",x"06",x"00",x"00"),
  1999 => (x"1e",x"3f",x"69",x"49"),
  2000 => (x"00",x"00",x"00",x"00"),
  2001 => (x"00",x"00",x"66",x"66"),
  2002 => (x"80",x"00",x"00",x"00"),
  2003 => (x"00",x"00",x"66",x"e6"),
  2004 => (x"08",x"08",x"00",x"00"),
  2005 => (x"22",x"22",x"14",x"14"),
  2006 => (x"14",x"14",x"00",x"00"),
  2007 => (x"14",x"14",x"14",x"14"),
  2008 => (x"22",x"22",x"00",x"00"),
  2009 => (x"08",x"08",x"14",x"14"),
  2010 => (x"03",x"02",x"00",x"00"),
  2011 => (x"06",x"0f",x"59",x"51"),
  2012 => (x"41",x"7f",x"3e",x"00"),
  2013 => (x"1e",x"1f",x"55",x"5d"),
  2014 => (x"7f",x"7e",x"00",x"00"),
  2015 => (x"7e",x"7f",x"09",x"09"),
  2016 => (x"7f",x"7f",x"00",x"00"),
  2017 => (x"36",x"7f",x"49",x"49"),
  2018 => (x"3e",x"1c",x"00",x"00"),
  2019 => (x"41",x"41",x"41",x"63"),
  2020 => (x"7f",x"7f",x"00",x"00"),
  2021 => (x"1c",x"3e",x"63",x"41"),
  2022 => (x"7f",x"7f",x"00",x"00"),
  2023 => (x"41",x"41",x"49",x"49"),
  2024 => (x"7f",x"7f",x"00",x"00"),
  2025 => (x"01",x"01",x"09",x"09"),
  2026 => (x"7f",x"3e",x"00",x"00"),
  2027 => (x"7a",x"7b",x"49",x"41"),
  2028 => (x"7f",x"7f",x"00",x"00"),
  2029 => (x"7f",x"7f",x"08",x"08"),
  2030 => (x"41",x"00",x"00",x"00"),
  2031 => (x"00",x"41",x"7f",x"7f"),
  2032 => (x"60",x"20",x"00",x"00"),
  2033 => (x"3f",x"7f",x"40",x"40"),
  2034 => (x"08",x"7f",x"7f",x"00"),
  2035 => (x"41",x"63",x"36",x"1c"),
  2036 => (x"7f",x"7f",x"00",x"00"),
  2037 => (x"40",x"40",x"40",x"40"),
  2038 => (x"06",x"7f",x"7f",x"00"),
  2039 => (x"7f",x"7f",x"06",x"0c"),
  2040 => (x"06",x"7f",x"7f",x"00"),
  2041 => (x"7f",x"7f",x"18",x"0c"),
  2042 => (x"7f",x"3e",x"00",x"00"),
  2043 => (x"3e",x"7f",x"41",x"41"),
  2044 => (x"7f",x"7f",x"00",x"00"),
  2045 => (x"06",x"0f",x"09",x"09"),
  2046 => (x"41",x"7f",x"3e",x"00"),
  2047 => (x"40",x"7e",x"7f",x"61"),
  2048 => (x"7f",x"7f",x"00",x"00"),
  2049 => (x"66",x"7f",x"19",x"09"),
  2050 => (x"6f",x"26",x"00",x"00"),
  2051 => (x"32",x"7b",x"59",x"4d"),
  2052 => (x"01",x"01",x"00",x"00"),
  2053 => (x"01",x"01",x"7f",x"7f"),
  2054 => (x"7f",x"3f",x"00",x"00"),
  2055 => (x"3f",x"7f",x"40",x"40"),
  2056 => (x"3f",x"0f",x"00",x"00"),
  2057 => (x"0f",x"3f",x"70",x"70"),
  2058 => (x"30",x"7f",x"7f",x"00"),
  2059 => (x"7f",x"7f",x"30",x"18"),
  2060 => (x"36",x"63",x"41",x"00"),
  2061 => (x"63",x"36",x"1c",x"1c"),
  2062 => (x"06",x"03",x"01",x"41"),
  2063 => (x"03",x"06",x"7c",x"7c"),
  2064 => (x"59",x"71",x"61",x"01"),
  2065 => (x"41",x"43",x"47",x"4d"),
  2066 => (x"7f",x"00",x"00",x"00"),
  2067 => (x"00",x"41",x"41",x"7f"),
  2068 => (x"06",x"03",x"01",x"00"),
  2069 => (x"60",x"30",x"18",x"0c"),
  2070 => (x"41",x"00",x"00",x"40"),
  2071 => (x"00",x"7f",x"7f",x"41"),
  2072 => (x"06",x"0c",x"08",x"00"),
  2073 => (x"08",x"0c",x"06",x"03"),
  2074 => (x"80",x"80",x"80",x"00"),
  2075 => (x"80",x"80",x"80",x"80"),
  2076 => (x"00",x"00",x"00",x"00"),
  2077 => (x"00",x"04",x"07",x"03"),
  2078 => (x"74",x"20",x"00",x"00"),
  2079 => (x"78",x"7c",x"54",x"54"),
  2080 => (x"7f",x"7f",x"00",x"00"),
  2081 => (x"38",x"7c",x"44",x"44"),
  2082 => (x"7c",x"38",x"00",x"00"),
  2083 => (x"00",x"44",x"44",x"44"),
  2084 => (x"7c",x"38",x"00",x"00"),
  2085 => (x"7f",x"7f",x"44",x"44"),
  2086 => (x"7c",x"38",x"00",x"00"),
  2087 => (x"18",x"5c",x"54",x"54"),
  2088 => (x"7e",x"04",x"00",x"00"),
  2089 => (x"00",x"05",x"05",x"7f"),
  2090 => (x"bc",x"18",x"00",x"00"),
  2091 => (x"7c",x"fc",x"a4",x"a4"),
  2092 => (x"7f",x"7f",x"00",x"00"),
  2093 => (x"78",x"7c",x"04",x"04"),
  2094 => (x"00",x"00",x"00",x"00"),
  2095 => (x"00",x"40",x"7d",x"3d"),
  2096 => (x"80",x"80",x"00",x"00"),
  2097 => (x"00",x"7d",x"fd",x"80"),
  2098 => (x"7f",x"7f",x"00",x"00"),
  2099 => (x"44",x"6c",x"38",x"10"),
  2100 => (x"00",x"00",x"00",x"00"),
  2101 => (x"00",x"40",x"7f",x"3f"),
  2102 => (x"0c",x"7c",x"7c",x"00"),
  2103 => (x"78",x"7c",x"0c",x"18"),
  2104 => (x"7c",x"7c",x"00",x"00"),
  2105 => (x"78",x"7c",x"04",x"04"),
  2106 => (x"7c",x"38",x"00",x"00"),
  2107 => (x"38",x"7c",x"44",x"44"),
  2108 => (x"fc",x"fc",x"00",x"00"),
  2109 => (x"18",x"3c",x"24",x"24"),
  2110 => (x"3c",x"18",x"00",x"00"),
  2111 => (x"fc",x"fc",x"24",x"24"),
  2112 => (x"7c",x"7c",x"00",x"00"),
  2113 => (x"08",x"0c",x"04",x"04"),
  2114 => (x"5c",x"48",x"00",x"00"),
  2115 => (x"20",x"74",x"54",x"54"),
  2116 => (x"3f",x"04",x"00",x"00"),
  2117 => (x"00",x"44",x"44",x"7f"),
  2118 => (x"7c",x"3c",x"00",x"00"),
  2119 => (x"7c",x"7c",x"40",x"40"),
  2120 => (x"3c",x"1c",x"00",x"00"),
  2121 => (x"1c",x"3c",x"60",x"60"),
  2122 => (x"60",x"7c",x"3c",x"00"),
  2123 => (x"3c",x"7c",x"60",x"30"),
  2124 => (x"38",x"6c",x"44",x"00"),
  2125 => (x"44",x"6c",x"38",x"10"),
  2126 => (x"bc",x"1c",x"00",x"00"),
  2127 => (x"1c",x"3c",x"60",x"e0"),
  2128 => (x"64",x"44",x"00",x"00"),
  2129 => (x"44",x"4c",x"5c",x"74"),
  2130 => (x"08",x"08",x"00",x"00"),
  2131 => (x"41",x"41",x"77",x"3e"),
  2132 => (x"00",x"00",x"00",x"00"),
  2133 => (x"00",x"00",x"7f",x"7f"),
  2134 => (x"41",x"41",x"00",x"00"),
  2135 => (x"08",x"08",x"3e",x"77"),
  2136 => (x"01",x"01",x"02",x"00"),
  2137 => (x"01",x"02",x"02",x"03"),
  2138 => (x"7f",x"7f",x"7f",x"00"),
  2139 => (x"7f",x"7f",x"7f",x"7f"),
  2140 => (x"1c",x"08",x"08",x"00"),
  2141 => (x"7f",x"3e",x"3e",x"1c"),
  2142 => (x"3e",x"7f",x"7f",x"7f"),
  2143 => (x"08",x"1c",x"1c",x"3e"),
  2144 => (x"18",x"10",x"00",x"08"),
  2145 => (x"10",x"18",x"7c",x"7c"),
  2146 => (x"30",x"10",x"00",x"00"),
  2147 => (x"10",x"30",x"7c",x"7c"),
  2148 => (x"60",x"30",x"10",x"00"),
  2149 => (x"06",x"1e",x"78",x"60"),
  2150 => (x"3c",x"66",x"42",x"00"),
  2151 => (x"42",x"66",x"3c",x"18"),
  2152 => (x"6a",x"38",x"78",x"00"),
  2153 => (x"38",x"6c",x"c6",x"c2"),
  2154 => (x"00",x"00",x"60",x"00"),
  2155 => (x"60",x"00",x"00",x"60"),
  2156 => (x"5b",x"5e",x"0e",x"00"),
  2157 => (x"1e",x"0e",x"5d",x"5c"),
  2158 => (x"f4",x"c2",x"4c",x"71"),
  2159 => (x"c0",x"4d",x"bf",x"fe"),
  2160 => (x"74",x"1e",x"c0",x"4b"),
  2161 => (x"87",x"c7",x"02",x"ab"),
  2162 => (x"c0",x"48",x"a6",x"c4"),
  2163 => (x"c4",x"87",x"c5",x"78"),
  2164 => (x"78",x"c1",x"48",x"a6"),
  2165 => (x"73",x"1e",x"66",x"c4"),
  2166 => (x"87",x"df",x"ee",x"49"),
  2167 => (x"e0",x"c0",x"86",x"c8"),
  2168 => (x"87",x"ef",x"ef",x"49"),
  2169 => (x"6a",x"4a",x"a5",x"c4"),
  2170 => (x"87",x"f0",x"f0",x"49"),
  2171 => (x"cb",x"87",x"c6",x"f1"),
  2172 => (x"c8",x"83",x"c1",x"85"),
  2173 => (x"ff",x"04",x"ab",x"b7"),
  2174 => (x"26",x"26",x"87",x"c7"),
  2175 => (x"26",x"4c",x"26",x"4d"),
  2176 => (x"1e",x"4f",x"26",x"4b"),
  2177 => (x"f5",x"c2",x"4a",x"71"),
  2178 => (x"f5",x"c2",x"5a",x"c2"),
  2179 => (x"78",x"c7",x"48",x"c2"),
  2180 => (x"87",x"dd",x"fe",x"49"),
  2181 => (x"73",x"1e",x"4f",x"26"),
  2182 => (x"c0",x"4a",x"71",x"1e"),
  2183 => (x"d3",x"03",x"aa",x"b7"),
  2184 => (x"e7",x"d5",x"c2",x"87"),
  2185 => (x"87",x"c4",x"05",x"bf"),
  2186 => (x"87",x"c2",x"4b",x"c1"),
  2187 => (x"d5",x"c2",x"4b",x"c0"),
  2188 => (x"87",x"c4",x"5b",x"eb"),
  2189 => (x"5a",x"eb",x"d5",x"c2"),
  2190 => (x"bf",x"e7",x"d5",x"c2"),
  2191 => (x"c1",x"9a",x"c1",x"4a"),
  2192 => (x"ec",x"49",x"a2",x"c0"),
  2193 => (x"48",x"fc",x"87",x"e8"),
  2194 => (x"bf",x"e7",x"d5",x"c2"),
  2195 => (x"87",x"ef",x"fe",x"78"),
  2196 => (x"c4",x"4a",x"71",x"1e"),
  2197 => (x"49",x"72",x"1e",x"66"),
  2198 => (x"26",x"87",x"fd",x"e9"),
  2199 => (x"c2",x"1e",x"4f",x"26"),
  2200 => (x"49",x"bf",x"e7",x"d5"),
  2201 => (x"c2",x"87",x"d7",x"e6"),
  2202 => (x"e8",x"48",x"f6",x"f4"),
  2203 => (x"f4",x"c2",x"78",x"bf"),
  2204 => (x"bf",x"ec",x"48",x"f2"),
  2205 => (x"f6",x"f4",x"c2",x"78"),
  2206 => (x"c3",x"49",x"4a",x"bf"),
  2207 => (x"b7",x"c8",x"99",x"ff"),
  2208 => (x"71",x"48",x"72",x"2a"),
  2209 => (x"fe",x"f4",x"c2",x"b0"),
  2210 => (x"0e",x"4f",x"26",x"58"),
  2211 => (x"5d",x"5c",x"5b",x"5e"),
  2212 => (x"ff",x"4b",x"71",x"0e"),
  2213 => (x"f4",x"c2",x"87",x"c8"),
  2214 => (x"50",x"c0",x"48",x"f1"),
  2215 => (x"fd",x"e5",x"49",x"73"),
  2216 => (x"4c",x"49",x"70",x"87"),
  2217 => (x"ee",x"cb",x"9c",x"c2"),
  2218 => (x"87",x"c3",x"cb",x"49"),
  2219 => (x"c2",x"4d",x"49",x"70"),
  2220 => (x"bf",x"97",x"f1",x"f4"),
  2221 => (x"87",x"e2",x"c1",x"05"),
  2222 => (x"c2",x"49",x"66",x"d0"),
  2223 => (x"99",x"bf",x"fa",x"f4"),
  2224 => (x"d4",x"87",x"d6",x"05"),
  2225 => (x"f4",x"c2",x"49",x"66"),
  2226 => (x"05",x"99",x"bf",x"f2"),
  2227 => (x"49",x"73",x"87",x"cb"),
  2228 => (x"70",x"87",x"cb",x"e5"),
  2229 => (x"c1",x"c1",x"02",x"98"),
  2230 => (x"fe",x"4c",x"c1",x"87"),
  2231 => (x"49",x"75",x"87",x"c0"),
  2232 => (x"70",x"87",x"d8",x"ca"),
  2233 => (x"87",x"c6",x"02",x"98"),
  2234 => (x"48",x"f1",x"f4",x"c2"),
  2235 => (x"f4",x"c2",x"50",x"c1"),
  2236 => (x"05",x"bf",x"97",x"f1"),
  2237 => (x"c2",x"87",x"e3",x"c0"),
  2238 => (x"49",x"bf",x"fa",x"f4"),
  2239 => (x"05",x"99",x"66",x"d0"),
  2240 => (x"c2",x"87",x"d6",x"ff"),
  2241 => (x"49",x"bf",x"f2",x"f4"),
  2242 => (x"05",x"99",x"66",x"d4"),
  2243 => (x"73",x"87",x"ca",x"ff"),
  2244 => (x"87",x"ca",x"e4",x"49"),
  2245 => (x"fe",x"05",x"98",x"70"),
  2246 => (x"48",x"74",x"87",x"ff"),
  2247 => (x"0e",x"87",x"dc",x"fb"),
  2248 => (x"5d",x"5c",x"5b",x"5e"),
  2249 => (x"c0",x"86",x"f4",x"0e"),
  2250 => (x"bf",x"ec",x"4c",x"4d"),
  2251 => (x"48",x"a6",x"c4",x"7e"),
  2252 => (x"bf",x"fe",x"f4",x"c2"),
  2253 => (x"c0",x"1e",x"c1",x"78"),
  2254 => (x"fd",x"49",x"c7",x"1e"),
  2255 => (x"86",x"c8",x"87",x"cd"),
  2256 => (x"cd",x"02",x"98",x"70"),
  2257 => (x"fb",x"49",x"ff",x"87"),
  2258 => (x"da",x"c1",x"87",x"cc"),
  2259 => (x"87",x"ce",x"e3",x"49"),
  2260 => (x"f4",x"c2",x"4d",x"c1"),
  2261 => (x"02",x"bf",x"97",x"f1"),
  2262 => (x"c3",x"d5",x"87",x"c3"),
  2263 => (x"f6",x"f4",x"c2",x"87"),
  2264 => (x"d5",x"c2",x"4b",x"bf"),
  2265 => (x"c0",x"05",x"bf",x"e7"),
  2266 => (x"fd",x"c3",x"87",x"e9"),
  2267 => (x"87",x"ee",x"e2",x"49"),
  2268 => (x"e2",x"49",x"fa",x"c3"),
  2269 => (x"49",x"73",x"87",x"e8"),
  2270 => (x"71",x"99",x"ff",x"c3"),
  2271 => (x"fb",x"49",x"c0",x"1e"),
  2272 => (x"49",x"73",x"87",x"ce"),
  2273 => (x"71",x"29",x"b7",x"c8"),
  2274 => (x"fb",x"49",x"c1",x"1e"),
  2275 => (x"86",x"c8",x"87",x"c2"),
  2276 => (x"c2",x"87",x"fa",x"c5"),
  2277 => (x"4b",x"bf",x"fa",x"f4"),
  2278 => (x"87",x"dd",x"02",x"9b"),
  2279 => (x"bf",x"e3",x"d5",x"c2"),
  2280 => (x"87",x"d7",x"c7",x"49"),
  2281 => (x"c4",x"05",x"98",x"70"),
  2282 => (x"d2",x"4b",x"c0",x"87"),
  2283 => (x"49",x"e0",x"c2",x"87"),
  2284 => (x"c2",x"87",x"fc",x"c6"),
  2285 => (x"c6",x"58",x"e7",x"d5"),
  2286 => (x"e3",x"d5",x"c2",x"87"),
  2287 => (x"73",x"78",x"c0",x"48"),
  2288 => (x"05",x"99",x"c2",x"49"),
  2289 => (x"eb",x"c3",x"87",x"cd"),
  2290 => (x"87",x"d2",x"e1",x"49"),
  2291 => (x"99",x"c2",x"49",x"70"),
  2292 => (x"fb",x"87",x"c2",x"02"),
  2293 => (x"c1",x"49",x"73",x"4c"),
  2294 => (x"87",x"cd",x"05",x"99"),
  2295 => (x"e0",x"49",x"f4",x"c3"),
  2296 => (x"49",x"70",x"87",x"fc"),
  2297 => (x"c2",x"02",x"99",x"c2"),
  2298 => (x"73",x"4c",x"fa",x"87"),
  2299 => (x"05",x"99",x"c8",x"49"),
  2300 => (x"f5",x"c3",x"87",x"cd"),
  2301 => (x"87",x"e6",x"e0",x"49"),
  2302 => (x"99",x"c2",x"49",x"70"),
  2303 => (x"c2",x"87",x"d4",x"02"),
  2304 => (x"02",x"bf",x"c2",x"f5"),
  2305 => (x"c1",x"48",x"87",x"c9"),
  2306 => (x"c6",x"f5",x"c2",x"88"),
  2307 => (x"ff",x"87",x"c2",x"58"),
  2308 => (x"73",x"4d",x"c1",x"4c"),
  2309 => (x"05",x"99",x"c4",x"49"),
  2310 => (x"f2",x"c3",x"87",x"ce"),
  2311 => (x"fd",x"df",x"ff",x"49"),
  2312 => (x"c2",x"49",x"70",x"87"),
  2313 => (x"87",x"db",x"02",x"99"),
  2314 => (x"bf",x"c2",x"f5",x"c2"),
  2315 => (x"b7",x"c7",x"48",x"7e"),
  2316 => (x"87",x"cb",x"03",x"a8"),
  2317 => (x"80",x"c1",x"48",x"6e"),
  2318 => (x"58",x"c6",x"f5",x"c2"),
  2319 => (x"fe",x"87",x"c2",x"c0"),
  2320 => (x"c3",x"4d",x"c1",x"4c"),
  2321 => (x"df",x"ff",x"49",x"fd"),
  2322 => (x"49",x"70",x"87",x"d4"),
  2323 => (x"d5",x"02",x"99",x"c2"),
  2324 => (x"c2",x"f5",x"c2",x"87"),
  2325 => (x"c9",x"c0",x"02",x"bf"),
  2326 => (x"c2",x"f5",x"c2",x"87"),
  2327 => (x"c0",x"78",x"c0",x"48"),
  2328 => (x"4c",x"fd",x"87",x"c2"),
  2329 => (x"fa",x"c3",x"4d",x"c1"),
  2330 => (x"f1",x"de",x"ff",x"49"),
  2331 => (x"c2",x"49",x"70",x"87"),
  2332 => (x"87",x"d9",x"02",x"99"),
  2333 => (x"bf",x"c2",x"f5",x"c2"),
  2334 => (x"a8",x"b7",x"c7",x"48"),
  2335 => (x"87",x"c9",x"c0",x"03"),
  2336 => (x"48",x"c2",x"f5",x"c2"),
  2337 => (x"c2",x"c0",x"78",x"c7"),
  2338 => (x"c1",x"4c",x"fc",x"87"),
  2339 => (x"ac",x"b7",x"c0",x"4d"),
  2340 => (x"87",x"d1",x"c0",x"03"),
  2341 => (x"c1",x"4a",x"66",x"c4"),
  2342 => (x"02",x"6a",x"82",x"d8"),
  2343 => (x"6a",x"87",x"c6",x"c0"),
  2344 => (x"73",x"49",x"74",x"4b"),
  2345 => (x"c3",x"1e",x"c0",x"0f"),
  2346 => (x"da",x"c1",x"1e",x"f0"),
  2347 => (x"87",x"db",x"f7",x"49"),
  2348 => (x"98",x"70",x"86",x"c8"),
  2349 => (x"87",x"e2",x"c0",x"02"),
  2350 => (x"c2",x"48",x"a6",x"c8"),
  2351 => (x"78",x"bf",x"c2",x"f5"),
  2352 => (x"cb",x"49",x"66",x"c8"),
  2353 => (x"48",x"66",x"c4",x"91"),
  2354 => (x"7e",x"70",x"80",x"71"),
  2355 => (x"c0",x"02",x"bf",x"6e"),
  2356 => (x"bf",x"6e",x"87",x"c8"),
  2357 => (x"49",x"66",x"c8",x"4b"),
  2358 => (x"9d",x"75",x"0f",x"73"),
  2359 => (x"87",x"c8",x"c0",x"02"),
  2360 => (x"bf",x"c2",x"f5",x"c2"),
  2361 => (x"87",x"c9",x"f3",x"49"),
  2362 => (x"bf",x"eb",x"d5",x"c2"),
  2363 => (x"87",x"dd",x"c0",x"02"),
  2364 => (x"87",x"c7",x"c2",x"49"),
  2365 => (x"c0",x"02",x"98",x"70"),
  2366 => (x"f5",x"c2",x"87",x"d3"),
  2367 => (x"f2",x"49",x"bf",x"c2"),
  2368 => (x"49",x"c0",x"87",x"ef"),
  2369 => (x"c2",x"87",x"cf",x"f4"),
  2370 => (x"c0",x"48",x"eb",x"d5"),
  2371 => (x"f3",x"8e",x"f4",x"78"),
  2372 => (x"5e",x"0e",x"87",x"e9"),
  2373 => (x"0e",x"5d",x"5c",x"5b"),
  2374 => (x"c2",x"4c",x"71",x"1e"),
  2375 => (x"49",x"bf",x"fe",x"f4"),
  2376 => (x"4d",x"a1",x"cd",x"c1"),
  2377 => (x"69",x"81",x"d1",x"c1"),
  2378 => (x"02",x"9c",x"74",x"7e"),
  2379 => (x"a5",x"c4",x"87",x"cf"),
  2380 => (x"c2",x"7b",x"74",x"4b"),
  2381 => (x"49",x"bf",x"fe",x"f4"),
  2382 => (x"6e",x"87",x"c8",x"f3"),
  2383 => (x"05",x"9c",x"74",x"7b"),
  2384 => (x"4b",x"c0",x"87",x"c4"),
  2385 => (x"4b",x"c1",x"87",x"c2"),
  2386 => (x"c9",x"f3",x"49",x"73"),
  2387 => (x"02",x"66",x"d4",x"87"),
  2388 => (x"da",x"49",x"87",x"c7"),
  2389 => (x"c2",x"4a",x"70",x"87"),
  2390 => (x"c2",x"4a",x"c0",x"87"),
  2391 => (x"26",x"5a",x"ef",x"d5"),
  2392 => (x"00",x"87",x"d8",x"f2"),
  2393 => (x"00",x"00",x"00",x"00"),
  2394 => (x"00",x"00",x"00",x"00"),
  2395 => (x"1e",x"00",x"00",x"00"),
  2396 => (x"c8",x"ff",x"4a",x"71"),
  2397 => (x"a1",x"72",x"49",x"bf"),
  2398 => (x"1e",x"4f",x"26",x"48"),
  2399 => (x"89",x"bf",x"c8",x"ff"),
  2400 => (x"c0",x"c0",x"c0",x"fe"),
  2401 => (x"01",x"a9",x"c0",x"c0"),
  2402 => (x"4a",x"c0",x"87",x"c4"),
  2403 => (x"4a",x"c1",x"87",x"c2"),
  2404 => (x"4f",x"26",x"48",x"72"),
  2405 => (x"5c",x"5b",x"5e",x"0e"),
  2406 => (x"4b",x"71",x"0e",x"5d"),
  2407 => (x"d0",x"4c",x"d4",x"ff"),
  2408 => (x"78",x"c0",x"48",x"66"),
  2409 => (x"db",x"ff",x"49",x"d6"),
  2410 => (x"ff",x"c3",x"87",x"f4"),
  2411 => (x"c3",x"49",x"6c",x"7c"),
  2412 => (x"4d",x"71",x"99",x"ff"),
  2413 => (x"99",x"f0",x"c3",x"49"),
  2414 => (x"05",x"a9",x"e0",x"c1"),
  2415 => (x"ff",x"c3",x"87",x"cb"),
  2416 => (x"c3",x"48",x"6c",x"7c"),
  2417 => (x"08",x"66",x"d0",x"98"),
  2418 => (x"7c",x"ff",x"c3",x"78"),
  2419 => (x"c8",x"49",x"4a",x"6c"),
  2420 => (x"7c",x"ff",x"c3",x"31"),
  2421 => (x"b2",x"71",x"4a",x"6c"),
  2422 => (x"31",x"c8",x"49",x"72"),
  2423 => (x"6c",x"7c",x"ff",x"c3"),
  2424 => (x"72",x"b2",x"71",x"4a"),
  2425 => (x"c3",x"31",x"c8",x"49"),
  2426 => (x"4a",x"6c",x"7c",x"ff"),
  2427 => (x"d0",x"ff",x"b2",x"71"),
  2428 => (x"78",x"e0",x"c0",x"48"),
  2429 => (x"c2",x"02",x"9b",x"73"),
  2430 => (x"75",x"7b",x"72",x"87"),
  2431 => (x"26",x"4d",x"26",x"48"),
  2432 => (x"26",x"4b",x"26",x"4c"),
  2433 => (x"4f",x"26",x"1e",x"4f"),
  2434 => (x"5c",x"5b",x"5e",x"0e"),
  2435 => (x"76",x"86",x"f8",x"0e"),
  2436 => (x"49",x"a6",x"c8",x"1e"),
  2437 => (x"c4",x"87",x"fd",x"fd"),
  2438 => (x"6e",x"4b",x"70",x"86"),
  2439 => (x"03",x"a8",x"c4",x"48"),
  2440 => (x"73",x"87",x"ca",x"c3"),
  2441 => (x"9a",x"f0",x"c3",x"4a"),
  2442 => (x"02",x"aa",x"d0",x"c1"),
  2443 => (x"e0",x"c1",x"87",x"c7"),
  2444 => (x"f8",x"c2",x"05",x"aa"),
  2445 => (x"c8",x"49",x"73",x"87"),
  2446 => (x"87",x"c3",x"02",x"99"),
  2447 => (x"73",x"87",x"c6",x"ff"),
  2448 => (x"c2",x"9c",x"c3",x"4c"),
  2449 => (x"cf",x"c1",x"05",x"ac"),
  2450 => (x"49",x"66",x"c4",x"87"),
  2451 => (x"1e",x"71",x"31",x"c9"),
  2452 => (x"c1",x"4a",x"66",x"c4"),
  2453 => (x"f5",x"c2",x"92",x"c8"),
  2454 => (x"81",x"72",x"49",x"c6"),
  2455 => (x"87",x"ef",x"d2",x"fe"),
  2456 => (x"1e",x"49",x"66",x"c4"),
  2457 => (x"ff",x"49",x"e3",x"c0"),
  2458 => (x"d8",x"87",x"d8",x"d9"),
  2459 => (x"ed",x"d8",x"ff",x"49"),
  2460 => (x"1e",x"c0",x"c8",x"87"),
  2461 => (x"49",x"f6",x"e3",x"c2"),
  2462 => (x"87",x"c4",x"eb",x"fd"),
  2463 => (x"c0",x"48",x"d0",x"ff"),
  2464 => (x"e3",x"c2",x"78",x"e0"),
  2465 => (x"66",x"d0",x"1e",x"f6"),
  2466 => (x"92",x"c8",x"c1",x"4a"),
  2467 => (x"49",x"c6",x"f5",x"c2"),
  2468 => (x"cd",x"fe",x"81",x"72"),
  2469 => (x"86",x"d0",x"87",x"f7"),
  2470 => (x"c1",x"05",x"ac",x"c1"),
  2471 => (x"66",x"c4",x"87",x"cf"),
  2472 => (x"71",x"31",x"c9",x"49"),
  2473 => (x"4a",x"66",x"c4",x"1e"),
  2474 => (x"c2",x"92",x"c8",x"c1"),
  2475 => (x"72",x"49",x"c6",x"f5"),
  2476 => (x"da",x"d1",x"fe",x"81"),
  2477 => (x"f6",x"e3",x"c2",x"87"),
  2478 => (x"4a",x"66",x"c8",x"1e"),
  2479 => (x"c2",x"92",x"c8",x"c1"),
  2480 => (x"72",x"49",x"c6",x"f5"),
  2481 => (x"c1",x"cc",x"fe",x"81"),
  2482 => (x"49",x"66",x"c8",x"87"),
  2483 => (x"49",x"e3",x"c0",x"1e"),
  2484 => (x"87",x"ef",x"d7",x"ff"),
  2485 => (x"d7",x"ff",x"49",x"d7"),
  2486 => (x"c0",x"c8",x"87",x"c4"),
  2487 => (x"f6",x"e3",x"c2",x"1e"),
  2488 => (x"c5",x"e9",x"fd",x"49"),
  2489 => (x"ff",x"86",x"d0",x"87"),
  2490 => (x"e0",x"c0",x"48",x"d0"),
  2491 => (x"fc",x"8e",x"f8",x"78"),
  2492 => (x"5e",x"0e",x"87",x"cd"),
  2493 => (x"0e",x"5d",x"5c",x"5b"),
  2494 => (x"ff",x"4d",x"71",x"1e"),
  2495 => (x"66",x"d4",x"4c",x"d4"),
  2496 => (x"b7",x"c3",x"48",x"7e"),
  2497 => (x"87",x"c5",x"06",x"a8"),
  2498 => (x"e3",x"c1",x"48",x"c0"),
  2499 => (x"fe",x"49",x"75",x"87"),
  2500 => (x"75",x"87",x"e3",x"e1"),
  2501 => (x"4b",x"66",x"c4",x"1e"),
  2502 => (x"c2",x"93",x"c8",x"c1"),
  2503 => (x"73",x"83",x"c6",x"f5"),
  2504 => (x"cf",x"c6",x"fe",x"49"),
  2505 => (x"6b",x"83",x"c8",x"87"),
  2506 => (x"48",x"d0",x"ff",x"4b"),
  2507 => (x"dd",x"78",x"e1",x"c8"),
  2508 => (x"c3",x"49",x"73",x"7c"),
  2509 => (x"7c",x"71",x"99",x"ff"),
  2510 => (x"b7",x"c8",x"49",x"73"),
  2511 => (x"99",x"ff",x"c3",x"29"),
  2512 => (x"49",x"73",x"7c",x"71"),
  2513 => (x"c3",x"29",x"b7",x"d0"),
  2514 => (x"7c",x"71",x"99",x"ff"),
  2515 => (x"b7",x"d8",x"49",x"73"),
  2516 => (x"c0",x"7c",x"71",x"29"),
  2517 => (x"7c",x"7c",x"7c",x"7c"),
  2518 => (x"7c",x"7c",x"7c",x"7c"),
  2519 => (x"7c",x"7c",x"7c",x"7c"),
  2520 => (x"c4",x"78",x"e0",x"c0"),
  2521 => (x"49",x"dc",x"1e",x"66"),
  2522 => (x"87",x"d7",x"d5",x"ff"),
  2523 => (x"48",x"73",x"86",x"c8"),
  2524 => (x"87",x"c9",x"fa",x"26"),
  2525 => (x"5c",x"5b",x"5e",x"0e"),
  2526 => (x"71",x"1e",x"0e",x"5d"),
  2527 => (x"4b",x"d4",x"ff",x"7e"),
  2528 => (x"f9",x"c2",x"1e",x"6e"),
  2529 => (x"c4",x"fe",x"49",x"e6"),
  2530 => (x"86",x"c4",x"87",x"ea"),
  2531 => (x"02",x"9d",x"4d",x"70"),
  2532 => (x"c2",x"87",x"c3",x"c3"),
  2533 => (x"4c",x"bf",x"ee",x"f9"),
  2534 => (x"df",x"fe",x"49",x"6e"),
  2535 => (x"d0",x"ff",x"87",x"d8"),
  2536 => (x"78",x"c5",x"c8",x"48"),
  2537 => (x"c0",x"7b",x"d6",x"c1"),
  2538 => (x"c1",x"7b",x"15",x"4a"),
  2539 => (x"b7",x"e0",x"c0",x"82"),
  2540 => (x"87",x"f5",x"04",x"aa"),
  2541 => (x"c4",x"48",x"d0",x"ff"),
  2542 => (x"78",x"c5",x"c8",x"78"),
  2543 => (x"c1",x"7b",x"d3",x"c1"),
  2544 => (x"74",x"78",x"c4",x"7b"),
  2545 => (x"fc",x"c1",x"02",x"9c"),
  2546 => (x"f6",x"e3",x"c2",x"87"),
  2547 => (x"4d",x"c0",x"c8",x"7e"),
  2548 => (x"ac",x"b7",x"c0",x"8c"),
  2549 => (x"c8",x"87",x"c6",x"03"),
  2550 => (x"c0",x"4d",x"a4",x"c0"),
  2551 => (x"e7",x"f0",x"c2",x"4c"),
  2552 => (x"d0",x"49",x"bf",x"97"),
  2553 => (x"87",x"d2",x"02",x"99"),
  2554 => (x"f9",x"c2",x"1e",x"c0"),
  2555 => (x"c7",x"fe",x"49",x"e6"),
  2556 => (x"86",x"c4",x"87",x"d8"),
  2557 => (x"c0",x"4a",x"49",x"70"),
  2558 => (x"e3",x"c2",x"87",x"ef"),
  2559 => (x"f9",x"c2",x"1e",x"f6"),
  2560 => (x"c7",x"fe",x"49",x"e6"),
  2561 => (x"86",x"c4",x"87",x"c4"),
  2562 => (x"ff",x"4a",x"49",x"70"),
  2563 => (x"c5",x"c8",x"48",x"d0"),
  2564 => (x"7b",x"d4",x"c1",x"78"),
  2565 => (x"7b",x"bf",x"97",x"6e"),
  2566 => (x"80",x"c1",x"48",x"6e"),
  2567 => (x"8d",x"c1",x"7e",x"70"),
  2568 => (x"87",x"f0",x"ff",x"05"),
  2569 => (x"c4",x"48",x"d0",x"ff"),
  2570 => (x"05",x"9a",x"72",x"78"),
  2571 => (x"48",x"c0",x"87",x"c5"),
  2572 => (x"c1",x"87",x"e5",x"c0"),
  2573 => (x"e6",x"f9",x"c2",x"1e"),
  2574 => (x"ec",x"c4",x"fe",x"49"),
  2575 => (x"74",x"86",x"c4",x"87"),
  2576 => (x"c4",x"fe",x"05",x"9c"),
  2577 => (x"48",x"d0",x"ff",x"87"),
  2578 => (x"c1",x"78",x"c5",x"c8"),
  2579 => (x"7b",x"c0",x"7b",x"d3"),
  2580 => (x"48",x"c1",x"78",x"c4"),
  2581 => (x"48",x"c0",x"87",x"c2"),
  2582 => (x"26",x"4d",x"26",x"26"),
  2583 => (x"26",x"4b",x"26",x"4c"),
  2584 => (x"5b",x"5e",x"0e",x"4f"),
  2585 => (x"4b",x"71",x"0e",x"5c"),
  2586 => (x"d8",x"02",x"66",x"cc"),
  2587 => (x"f0",x"c0",x"4c",x"87"),
  2588 => (x"87",x"d8",x"02",x"8c"),
  2589 => (x"8a",x"c1",x"4a",x"74"),
  2590 => (x"8a",x"87",x"d1",x"02"),
  2591 => (x"8a",x"87",x"cd",x"02"),
  2592 => (x"d7",x"87",x"c9",x"02"),
  2593 => (x"fb",x"49",x"73",x"87"),
  2594 => (x"87",x"d0",x"87",x"ea"),
  2595 => (x"49",x"c0",x"1e",x"74"),
  2596 => (x"74",x"87",x"df",x"f9"),
  2597 => (x"f9",x"49",x"73",x"1e"),
  2598 => (x"86",x"c8",x"87",x"d8"),
  2599 => (x"00",x"87",x"fc",x"fe"),
  2600 => (x"c9",x"e3",x"c2",x"1e"),
  2601 => (x"b9",x"c1",x"49",x"bf"),
  2602 => (x"59",x"cd",x"e3",x"c2"),
  2603 => (x"c3",x"48",x"d4",x"ff"),
  2604 => (x"d0",x"ff",x"78",x"ff"),
  2605 => (x"78",x"e1",x"c8",x"48"),
  2606 => (x"c1",x"48",x"d4",x"ff"),
  2607 => (x"71",x"31",x"c4",x"78"),
  2608 => (x"48",x"d0",x"ff",x"78"),
  2609 => (x"26",x"78",x"e0",x"c0"),
  2610 => (x"00",x"00",x"00",x"4f"),
  2611 => (x"00",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

