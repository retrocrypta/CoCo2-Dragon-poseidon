library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"f0fac287",
    12 => x"86c0c64e",
    13 => x"49f0fac2",
    14 => x"48d0e3c2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087dbe3",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"4a66c41e",
    47 => x"51124871",
    48 => x"2687fb05",
    49 => x"1e731e4f",
    50 => x"c0029a72",
    51 => x"48c087e7",
    52 => x"a9724bc1",
    53 => x"7287d106",
    54 => x"87c90682",
    55 => x"a9728373",
    56 => x"c387f401",
    57 => x"3ab2c187",
    58 => x"8903a972",
    59 => x"c1078073",
    60 => x"f3052b2a",
    61 => x"264b2687",
    62 => x"1e751e4f",
    63 => x"b7714dc4",
    64 => x"b9ff04a1",
    65 => x"bdc381c1",
    66 => x"a2b77207",
    67 => x"c1baff04",
    68 => x"07bdc182",
    69 => x"c187eefe",
    70 => x"b8ff042d",
    71 => x"2d0780c1",
    72 => x"c1b9ff04",
    73 => x"4d260781",
    74 => x"111e4f26",
    75 => x"08d4ff48",
    76 => x"4866c478",
    77 => x"a6c888c1",
    78 => x"05987058",
    79 => x"4f2687ed",
    80 => x"48d4ff1e",
    81 => x"6878ffc3",
    82 => x"4866c451",
    83 => x"a6c888c1",
    84 => x"05987058",
    85 => x"4f2687eb",
    86 => x"ff1e731e",
    87 => x"ffc34bd4",
    88 => x"c34a6b7b",
    89 => x"496b7bff",
    90 => x"b17232c8",
    91 => x"6b7bffc3",
    92 => x"7131c84a",
    93 => x"7bffc3b2",
    94 => x"32c8496b",
    95 => x"4871b172",
    96 => x"4d2687c4",
    97 => x"4b264c26",
    98 => x"5e0e4f26",
    99 => x"0e5d5c5b",
   100 => x"d4ff4a71",
   101 => x"c349724c",
   102 => x"7c7199ff",
   103 => x"bfd0e3c2",
   104 => x"d087c805",
   105 => x"30c94866",
   106 => x"d058a6d4",
   107 => x"29d84966",
   108 => x"7199ffc3",
   109 => x"4966d07c",
   110 => x"ffc329d0",
   111 => x"d07c7199",
   112 => x"29c84966",
   113 => x"7199ffc3",
   114 => x"4966d07c",
   115 => x"7199ffc3",
   116 => x"d049727c",
   117 => x"99ffc329",
   118 => x"4b6c7c71",
   119 => x"4dfff0c9",
   120 => x"05abffc3",
   121 => x"ffc387d0",
   122 => x"c14b6c7c",
   123 => x"87c6028d",
   124 => x"02abffc3",
   125 => x"487387f0",
   126 => x"1e87c7fe",
   127 => x"d4ff49c0",
   128 => x"78ffc348",
   129 => x"c8c381c1",
   130 => x"f104a9b7",
   131 => x"1e4f2687",
   132 => x"87e71e73",
   133 => x"4bdff8c4",
   134 => x"ffc01ec0",
   135 => x"49f7c1f0",
   136 => x"c487e7fd",
   137 => x"05a8c186",
   138 => x"ff87eac0",
   139 => x"ffc348d4",
   140 => x"c0c0c178",
   141 => x"1ec0c0c0",
   142 => x"c1f0e1c0",
   143 => x"c9fd49e9",
   144 => x"7086c487",
   145 => x"87ca0598",
   146 => x"c348d4ff",
   147 => x"48c178ff",
   148 => x"e6fe87cb",
   149 => x"058bc187",
   150 => x"c087fdfe",
   151 => x"87e6fc48",
   152 => x"ff1e731e",
   153 => x"ffc348d4",
   154 => x"c04bd378",
   155 => x"f0ffc01e",
   156 => x"fc49c1c1",
   157 => x"86c487d4",
   158 => x"ca059870",
   159 => x"48d4ff87",
   160 => x"c178ffc3",
   161 => x"fd87cb48",
   162 => x"8bc187f1",
   163 => x"87dbff05",
   164 => x"f1fb48c0",
   165 => x"5b5e0e87",
   166 => x"d4ff0e5c",
   167 => x"87dbfd4c",
   168 => x"c01eeac6",
   169 => x"c8c1f0e1",
   170 => x"87defb49",
   171 => x"a8c186c4",
   172 => x"fe87c802",
   173 => x"48c087ea",
   174 => x"fa87e2c1",
   175 => x"497087da",
   176 => x"99ffffcf",
   177 => x"02a9eac6",
   178 => x"d3fe87c8",
   179 => x"c148c087",
   180 => x"ffc387cb",
   181 => x"4bf1c07c",
   182 => x"7087f4fc",
   183 => x"ebc00298",
   184 => x"c01ec087",
   185 => x"fac1f0ff",
   186 => x"87defa49",
   187 => x"987086c4",
   188 => x"c387d905",
   189 => x"496c7cff",
   190 => x"7c7cffc3",
   191 => x"c0c17c7c",
   192 => x"87c40299",
   193 => x"87d548c1",
   194 => x"87d148c0",
   195 => x"c405abc2",
   196 => x"c848c087",
   197 => x"058bc187",
   198 => x"c087fdfe",
   199 => x"87e4f948",
   200 => x"c21e731e",
   201 => x"c148d0e3",
   202 => x"ff4bc778",
   203 => x"78c248d0",
   204 => x"ff87c8fb",
   205 => x"78c348d0",
   206 => x"e5c01ec0",
   207 => x"49c0c1d0",
   208 => x"c487c7f9",
   209 => x"05a8c186",
   210 => x"c24b87c1",
   211 => x"87c505ab",
   212 => x"f9c048c0",
   213 => x"058bc187",
   214 => x"fc87d0ff",
   215 => x"e3c287f7",
   216 => x"987058d4",
   217 => x"c187cd05",
   218 => x"f0ffc01e",
   219 => x"f849d0c1",
   220 => x"86c487d8",
   221 => x"c348d4ff",
   222 => x"e0c478ff",
   223 => x"d8e3c287",
   224 => x"48d0ff58",
   225 => x"d4ff78c2",
   226 => x"78ffc348",
   227 => x"f5f748c1",
   228 => x"5b5e0e87",
   229 => x"710e5d5c",
   230 => x"4dffc34a",
   231 => x"754cd4ff",
   232 => x"48d0ff7c",
   233 => x"7578c3c4",
   234 => x"c01e727c",
   235 => x"d8c1f0ff",
   236 => x"87d6f749",
   237 => x"987086c4",
   238 => x"c087c502",
   239 => x"87f0c048",
   240 => x"fec37c75",
   241 => x"1ec0c87c",
   242 => x"f54966d4",
   243 => x"86c487dc",
   244 => x"7c757c75",
   245 => x"dad87c75",
   246 => x"7c754be0",
   247 => x"0599496c",
   248 => x"8bc187c5",
   249 => x"7587f305",
   250 => x"48d0ff7c",
   251 => x"48c178c2",
   252 => x"1e87cff6",
   253 => x"ff4ad4ff",
   254 => x"d1c448d0",
   255 => x"7affc378",
   256 => x"f80589c1",
   257 => x"1e4f2687",
   258 => x"4b711e73",
   259 => x"dfcdeec5",
   260 => x"48d4ff4a",
   261 => x"6878ffc3",
   262 => x"a8fec348",
   263 => x"c187c502",
   264 => x"87ed058a",
   265 => x"c5059a72",
   266 => x"c048c087",
   267 => x"9b7387ea",
   268 => x"c887cc02",
   269 => x"49731e66",
   270 => x"c487c5f4",
   271 => x"c887c686",
   272 => x"eefe4966",
   273 => x"48d4ff87",
   274 => x"7878ffc3",
   275 => x"c5059b73",
   276 => x"48d0ff87",
   277 => x"48c178d0",
   278 => x"1e87ebf4",
   279 => x"4a711e73",
   280 => x"d4ff4bc0",
   281 => x"78ffc348",
   282 => x"c448d0ff",
   283 => x"d4ff78c3",
   284 => x"78ffc348",
   285 => x"ffc01e72",
   286 => x"49d1c1f0",
   287 => x"c487cbf4",
   288 => x"05987086",
   289 => x"c0c887cd",
   290 => x"4966cc1e",
   291 => x"c487f8fd",
   292 => x"ff4b7086",
   293 => x"78c248d0",
   294 => x"e9f34873",
   295 => x"5b5e0e87",
   296 => x"c00e5d5c",
   297 => x"f0ffc01e",
   298 => x"f349c9c1",
   299 => x"1ed287dc",
   300 => x"49d8e3c2",
   301 => x"c887d0fd",
   302 => x"c14cc086",
   303 => x"acb7d284",
   304 => x"c287f804",
   305 => x"bf97d8e3",
   306 => x"99c0c349",
   307 => x"05a9c0c1",
   308 => x"c287e7c0",
   309 => x"bf97dfe3",
   310 => x"c231d049",
   311 => x"bf97e0e3",
   312 => x"7232c84a",
   313 => x"e1e3c2b1",
   314 => x"b14abf97",
   315 => x"ffcf4c71",
   316 => x"c19cffff",
   317 => x"c134ca84",
   318 => x"e3c287e7",
   319 => x"49bf97e1",
   320 => x"99c631c1",
   321 => x"97e2e3c2",
   322 => x"b7c74abf",
   323 => x"c2b1722a",
   324 => x"bf97dde3",
   325 => x"9dcf4d4a",
   326 => x"97dee3c2",
   327 => x"9ac34abf",
   328 => x"e3c232ca",
   329 => x"4bbf97df",
   330 => x"b27333c2",
   331 => x"97e0e3c2",
   332 => x"c0c34bbf",
   333 => x"2bb7c69b",
   334 => x"81c2b273",
   335 => x"307148c1",
   336 => x"48c14970",
   337 => x"4d703075",
   338 => x"84c14c72",
   339 => x"c0c89471",
   340 => x"cc06adb7",
   341 => x"b734c187",
   342 => x"b7c0c82d",
   343 => x"f4ff01ad",
   344 => x"f0487487",
   345 => x"5e0e87dc",
   346 => x"0e5d5c5b",
   347 => x"ebc286f8",
   348 => x"78c048fe",
   349 => x"1ef6e3c2",
   350 => x"defb49c0",
   351 => x"7086c487",
   352 => x"87c50598",
   353 => x"cec948c0",
   354 => x"c14dc087",
   355 => x"c1fac07e",
   356 => x"e4c249bf",
   357 => x"c8714aec",
   358 => x"87ceeb4b",
   359 => x"c2059870",
   360 => x"c07ec087",
   361 => x"49bffdf9",
   362 => x"4ac8e5c2",
   363 => x"ea4bc871",
   364 => x"987087f8",
   365 => x"c087c205",
   366 => x"c0026e7e",
   367 => x"eac287fd",
   368 => x"c24dbffc",
   369 => x"bf9ff4eb",
   370 => x"d6c5487e",
   371 => x"c705a8ea",
   372 => x"fceac287",
   373 => x"87ce4dbf",
   374 => x"e9ca486e",
   375 => x"c502a8d5",
   376 => x"c748c087",
   377 => x"e3c287f1",
   378 => x"49751ef6",
   379 => x"c487ecf9",
   380 => x"05987086",
   381 => x"48c087c5",
   382 => x"c087dcc7",
   383 => x"49bffdf9",
   384 => x"4ac8e5c2",
   385 => x"e94bc871",
   386 => x"987087e0",
   387 => x"c287c805",
   388 => x"c148feeb",
   389 => x"c087da78",
   390 => x"49bfc1fa",
   391 => x"4aece4c2",
   392 => x"e94bc871",
   393 => x"987087c4",
   394 => x"87c5c002",
   395 => x"e6c648c0",
   396 => x"f4ebc287",
   397 => x"c149bf97",
   398 => x"c005a9d5",
   399 => x"ebc287cd",
   400 => x"49bf97f5",
   401 => x"02a9eac2",
   402 => x"c087c5c0",
   403 => x"87c7c648",
   404 => x"97f6e3c2",
   405 => x"c3487ebf",
   406 => x"c002a8e9",
   407 => x"486e87ce",
   408 => x"02a8ebc3",
   409 => x"c087c5c0",
   410 => x"87ebc548",
   411 => x"97c1e4c2",
   412 => x"059949bf",
   413 => x"c287ccc0",
   414 => x"bf97c2e4",
   415 => x"02a9c249",
   416 => x"c087c5c0",
   417 => x"87cfc548",
   418 => x"97c3e4c2",
   419 => x"ebc248bf",
   420 => x"4c7058fa",
   421 => x"c288c148",
   422 => x"c258feeb",
   423 => x"bf97c4e4",
   424 => x"c2817549",
   425 => x"bf97c5e4",
   426 => x"7232c84a",
   427 => x"f0c27ea1",
   428 => x"786e48cb",
   429 => x"97c6e4c2",
   430 => x"a6c848bf",
   431 => x"feebc258",
   432 => x"d4c202bf",
   433 => x"fdf9c087",
   434 => x"e5c249bf",
   435 => x"c8714ac8",
   436 => x"87d6e64b",
   437 => x"c0029870",
   438 => x"48c087c5",
   439 => x"c287f8c3",
   440 => x"4cbff6eb",
   441 => x"5cdff0c2",
   442 => x"97dbe4c2",
   443 => x"31c849bf",
   444 => x"97dae4c2",
   445 => x"49a14abf",
   446 => x"97dce4c2",
   447 => x"32d04abf",
   448 => x"c249a172",
   449 => x"bf97dde4",
   450 => x"7232d84a",
   451 => x"66c449a1",
   452 => x"cbf0c291",
   453 => x"f0c281bf",
   454 => x"e4c259d3",
   455 => x"4abf97e3",
   456 => x"e4c232c8",
   457 => x"4bbf97e2",
   458 => x"e4c24aa2",
   459 => x"4bbf97e4",
   460 => x"a27333d0",
   461 => x"e5e4c24a",
   462 => x"cf4bbf97",
   463 => x"7333d89b",
   464 => x"f0c24aa2",
   465 => x"f0c25ad7",
   466 => x"c24abfd3",
   467 => x"c292748a",
   468 => x"7248d7f0",
   469 => x"cac178a1",
   470 => x"c8e4c287",
   471 => x"c849bf97",
   472 => x"c7e4c231",
   473 => x"a14abf97",
   474 => x"c6ecc249",
   475 => x"c2ecc259",
   476 => x"31c549bf",
   477 => x"c981ffc7",
   478 => x"dff0c229",
   479 => x"cde4c259",
   480 => x"c84abf97",
   481 => x"cce4c232",
   482 => x"a24bbf97",
   483 => x"9266c44a",
   484 => x"f0c2826e",
   485 => x"f0c25adb",
   486 => x"78c048d3",
   487 => x"48cff0c2",
   488 => x"c278a172",
   489 => x"c248dff0",
   490 => x"78bfd3f0",
   491 => x"48e3f0c2",
   492 => x"bfd7f0c2",
   493 => x"feebc278",
   494 => x"c9c002bf",
   495 => x"c4487487",
   496 => x"c07e7030",
   497 => x"f0c287c9",
   498 => x"c448bfdb",
   499 => x"c27e7030",
   500 => x"6e48c2ec",
   501 => x"f848c178",
   502 => x"264d268e",
   503 => x"264b264c",
   504 => x"5b5e0e4f",
   505 => x"710e5d5c",
   506 => x"feebc24a",
   507 => x"87cb02bf",
   508 => x"2bc74b72",
   509 => x"ffc14c72",
   510 => x"7287c99c",
   511 => x"722bc84b",
   512 => x"9cffc34c",
   513 => x"bfcbf0c2",
   514 => x"f9f9c083",
   515 => x"d902abbf",
   516 => x"fdf9c087",
   517 => x"f6e3c25b",
   518 => x"f049731e",
   519 => x"86c487fd",
   520 => x"c5059870",
   521 => x"c048c087",
   522 => x"ebc287e6",
   523 => x"d202bffe",
   524 => x"c4497487",
   525 => x"f6e3c291",
   526 => x"cf4d6981",
   527 => x"ffffffff",
   528 => x"7487cb9d",
   529 => x"c291c249",
   530 => x"9f81f6e3",
   531 => x"48754d69",
   532 => x"0e87c6fe",
   533 => x"5d5c5b5e",
   534 => x"4d711e0e",
   535 => x"49c11ec0",
   536 => x"c487fed0",
   537 => x"9c4c7086",
   538 => x"87c2c102",
   539 => x"4ac6ecc2",
   540 => x"dfff4975",
   541 => x"987087d9",
   542 => x"87f2c002",
   543 => x"49754a74",
   544 => x"dfff4bcb",
   545 => x"987087fe",
   546 => x"87e2c002",
   547 => x"9c741ec0",
   548 => x"c487c702",
   549 => x"78c048a6",
   550 => x"a6c487c5",
   551 => x"c478c148",
   552 => x"fccf4966",
   553 => x"7086c487",
   554 => x"fe059c4c",
   555 => x"487487fe",
   556 => x"87e5fc26",
   557 => x"5c5b5e0e",
   558 => x"86f80e5d",
   559 => x"059b4b71",
   560 => x"48c087c5",
   561 => x"c887ddc2",
   562 => x"7dc04da3",
   563 => x"c70266d8",
   564 => x"9766d887",
   565 => x"87c505bf",
   566 => x"c7c248c0",
   567 => x"4966d887",
   568 => x"7087f0fd",
   569 => x"c1026e7e",
   570 => x"496e87f8",
   571 => x"7d6981dc",
   572 => x"81da496e",
   573 => x"9f4ca3c4",
   574 => x"ebc27c69",
   575 => x"d002bffe",
   576 => x"d4496e87",
   577 => x"49699f81",
   578 => x"ffffc04a",
   579 => x"c232d09a",
   580 => x"724ac087",
   581 => x"806c4849",
   582 => x"7bc07c70",
   583 => x"6c49a3cc",
   584 => x"49a3d079",
   585 => x"a6c479c0",
   586 => x"d478c048",
   587 => x"66c44aa3",
   588 => x"7291c849",
   589 => x"41c049a1",
   590 => x"66c4796c",
   591 => x"c880c148",
   592 => x"b7c658a6",
   593 => x"e2ff04a8",
   594 => x"c94a6d87",
   595 => x"c049722a",
   596 => x"ddff4af0",
   597 => x"4a7087ef",
   598 => x"49a3c4c1",
   599 => x"486e7972",
   600 => x"48c087c2",
   601 => x"f0f98ef8",
   602 => x"5b5e0e87",
   603 => x"710e5d5c",
   604 => x"f9f9c04c",
   605 => x"7478ff48",
   606 => x"cac1029c",
   607 => x"49a4c887",
   608 => x"c2c10269",
   609 => x"4a66d087",
   610 => x"d482496c",
   611 => x"66d05aa6",
   612 => x"ebc2b94d",
   613 => x"ff4abffa",
   614 => x"719972ba",
   615 => x"e4c00299",
   616 => x"4ba4c487",
   617 => x"f8f8496b",
   618 => x"c27b7087",
   619 => x"49bff6eb",
   620 => x"7c71816c",
   621 => x"ebc2b975",
   622 => x"ff4abffa",
   623 => x"719972ba",
   624 => x"dcff0599",
   625 => x"f87c7587",
   626 => x"731e87cf",
   627 => x"9b4b711e",
   628 => x"c887c702",
   629 => x"056949a3",
   630 => x"48c087c5",
   631 => x"c287ebc0",
   632 => x"4abfcff0",
   633 => x"6949a3c4",
   634 => x"c289c249",
   635 => x"91bff6eb",
   636 => x"c24aa271",
   637 => x"49bffaeb",
   638 => x"a271996b",
   639 => x"1e66c84a",
   640 => x"d6e94972",
   641 => x"7086c487",
   642 => x"d0f74849",
   643 => x"1e731e87",
   644 => x"029b4b71",
   645 => x"a3c887c7",
   646 => x"c5056949",
   647 => x"c048c087",
   648 => x"f0c287eb",
   649 => x"c44abfcf",
   650 => x"496949a3",
   651 => x"ebc289c2",
   652 => x"7191bff6",
   653 => x"ebc24aa2",
   654 => x"6b49bffa",
   655 => x"4aa27199",
   656 => x"721e66c8",
   657 => x"87c9e549",
   658 => x"497086c4",
   659 => x"87cdf648",
   660 => x"5c5b5e0e",
   661 => x"86f80e5d",
   662 => x"a6c44b71",
   663 => x"c878ff48",
   664 => x"4d6949a3",
   665 => x"a3d44cc0",
   666 => x"c849744a",
   667 => x"49a17291",
   668 => x"66d84969",
   669 => x"70887148",
   670 => x"a966d87e",
   671 => x"6e87ca01",
   672 => x"87c506ad",
   673 => x"6e5ca6c8",
   674 => x"c684c14d",
   675 => x"ff04acb7",
   676 => x"66c487d4",
   677 => x"f48ef848",
   678 => x"5e0e87ff",
   679 => x"0e5d5c5b",
   680 => x"a6c886ec",
   681 => x"48a6c859",
   682 => x"ffffffc1",
   683 => x"c478ffff",
   684 => x"c078ff80",
   685 => x"c44cc04d",
   686 => x"83d44b66",
   687 => x"91c84974",
   688 => x"7549a173",
   689 => x"7392c84a",
   690 => x"49697ea2",
   691 => x"d489bf6e",
   692 => x"ad7459a6",
   693 => x"d087c605",
   694 => x"bf6e48a6",
   695 => x"4866d078",
   696 => x"04a8b7c0",
   697 => x"66d087cf",
   698 => x"a966c849",
   699 => x"d087c603",
   700 => x"a6cc5ca6",
   701 => x"c684c159",
   702 => x"fe04acb7",
   703 => x"85c187f9",
   704 => x"04adb7c6",
   705 => x"cc87eefe",
   706 => x"8eec4866",
   707 => x"0e87caf3",
   708 => x"5d5c5b5e",
   709 => x"7186f00e",
   710 => x"66e0c04b",
   711 => x"732cc94c",
   712 => x"e1c3029b",
   713 => x"49a3c887",
   714 => x"d9c30269",
   715 => x"49a3d087",
   716 => x"7966e0c0",
   717 => x"02ac7e6b",
   718 => x"c287cbc3",
   719 => x"49bffaeb",
   720 => x"4a71b9ff",
   721 => x"48719a74",
   722 => x"a6cc986e",
   723 => x"4da3c458",
   724 => x"6d48a6c4",
   725 => x"aa66c878",
   726 => x"7487c505",
   727 => x"87d1c27b",
   728 => x"49731e72",
   729 => x"c487e9fb",
   730 => x"487e7086",
   731 => x"04a8b7c0",
   732 => x"a3d487d0",
   733 => x"c8496e4a",
   734 => x"49a17291",
   735 => x"7d697b21",
   736 => x"7bc087c7",
   737 => x"6949a3cc",
   738 => x"1e66c87d",
   739 => x"fffa4973",
   740 => x"7086c487",
   741 => x"a3c4c17e",
   742 => x"48a6cc49",
   743 => x"66c87869",
   744 => x"a866cc48",
   745 => x"6e87c906",
   746 => x"a8b7c048",
   747 => x"87e0c004",
   748 => x"b7c0486e",
   749 => x"ecc004a8",
   750 => x"4aa3d487",
   751 => x"91c8496e",
   752 => x"c849a172",
   753 => x"88694866",
   754 => x"66cc4970",
   755 => x"87d506a9",
   756 => x"c5fb4973",
   757 => x"d4497087",
   758 => x"91c84aa3",
   759 => x"c849a172",
   760 => x"66c44166",
   761 => x"748c6b79",
   762 => x"49731e49",
   763 => x"c487faf5",
   764 => x"66e0c086",
   765 => x"99ffc749",
   766 => x"c287cb02",
   767 => x"731ef6e3",
   768 => x"87c6f749",
   769 => x"8ef086c4",
   770 => x"1e87ceef",
   771 => x"4b711e73",
   772 => x"e4c0029b",
   773 => x"e3f0c287",
   774 => x"c24a735b",
   775 => x"f6ebc28a",
   776 => x"c29249bf",
   777 => x"48bfcff0",
   778 => x"f0c28072",
   779 => x"487158e7",
   780 => x"ecc230c4",
   781 => x"edc058c6",
   782 => x"dff0c287",
   783 => x"d3f0c248",
   784 => x"f0c278bf",
   785 => x"f0c248e3",
   786 => x"c278bfd7",
   787 => x"02bffeeb",
   788 => x"ebc287c9",
   789 => x"c449bff6",
   790 => x"c287c731",
   791 => x"49bfdbf0",
   792 => x"ecc231c4",
   793 => x"f4ed59c6",
   794 => x"5b5e0e87",
   795 => x"4a710e5c",
   796 => x"9a724bc0",
   797 => x"87e1c002",
   798 => x"9f49a2da",
   799 => x"ebc24b69",
   800 => x"cf02bffe",
   801 => x"49a2d487",
   802 => x"4c49699f",
   803 => x"9cffffc0",
   804 => x"87c234d0",
   805 => x"49744cc0",
   806 => x"fd4973b3",
   807 => x"faec87ed",
   808 => x"5b5e0e87",
   809 => x"f40e5d5c",
   810 => x"c04a7186",
   811 => x"029a727e",
   812 => x"e3c287d8",
   813 => x"78c048f2",
   814 => x"48eae3c2",
   815 => x"bfe3f0c2",
   816 => x"eee3c278",
   817 => x"dff0c248",
   818 => x"ecc278bf",
   819 => x"50c048d3",
   820 => x"bfc2ecc2",
   821 => x"f2e3c249",
   822 => x"aa714abf",
   823 => x"87c0c403",
   824 => x"99cf4972",
   825 => x"87e1c005",
   826 => x"1ef6e3c2",
   827 => x"bfeae3c2",
   828 => x"eae3c249",
   829 => x"78a1c148",
   830 => x"deddff71",
   831 => x"c086c487",
   832 => x"c248f5f9",
   833 => x"cc78f6e3",
   834 => x"f5f9c087",
   835 => x"e0c048bf",
   836 => x"f9f9c080",
   837 => x"f2e3c258",
   838 => x"80c148bf",
   839 => x"58f6e3c2",
   840 => x"000e7527",
   841 => x"bf97bf00",
   842 => x"c2029d4d",
   843 => x"e5c387e2",
   844 => x"dbc202ad",
   845 => x"f5f9c087",
   846 => x"a3cb4bbf",
   847 => x"cf4c1149",
   848 => x"d2c105ac",
   849 => x"df497587",
   850 => x"cd89c199",
   851 => x"c6ecc291",
   852 => x"4aa3c181",
   853 => x"a3c35112",
   854 => x"c551124a",
   855 => x"51124aa3",
   856 => x"124aa3c7",
   857 => x"4aa3c951",
   858 => x"a3ce5112",
   859 => x"d051124a",
   860 => x"51124aa3",
   861 => x"124aa3d2",
   862 => x"4aa3d451",
   863 => x"a3d65112",
   864 => x"d851124a",
   865 => x"51124aa3",
   866 => x"124aa3dc",
   867 => x"4aa3de51",
   868 => x"7ec15112",
   869 => x"7487f9c0",
   870 => x"0599c849",
   871 => x"7487eac0",
   872 => x"0599d049",
   873 => x"66dc87d0",
   874 => x"87cac002",
   875 => x"66dc4973",
   876 => x"0298700f",
   877 => x"056e87d3",
   878 => x"c287c6c0",
   879 => x"c048c6ec",
   880 => x"f5f9c050",
   881 => x"e7c248bf",
   882 => x"d3ecc287",
   883 => x"7e50c048",
   884 => x"bfc2ecc2",
   885 => x"f2e3c249",
   886 => x"aa714abf",
   887 => x"87c0fc04",
   888 => x"bfe3f0c2",
   889 => x"87c8c005",
   890 => x"bffeebc2",
   891 => x"87fec102",
   892 => x"48f9f9c0",
   893 => x"e3c278ff",
   894 => x"e749bfee",
   895 => x"497087e3",
   896 => x"59f2e3c2",
   897 => x"c248a6c4",
   898 => x"78bfeee3",
   899 => x"bffeebc2",
   900 => x"87d8c002",
   901 => x"cf4966c4",
   902 => x"f8ffffff",
   903 => x"c002a999",
   904 => x"4dc087c5",
   905 => x"c187e1c0",
   906 => x"87dcc04d",
   907 => x"cf4966c4",
   908 => x"a999f8ff",
   909 => x"87c8c002",
   910 => x"c048a6c8",
   911 => x"87c5c078",
   912 => x"c148a6c8",
   913 => x"4d66c878",
   914 => x"c0059d75",
   915 => x"66c487e0",
   916 => x"c289c249",
   917 => x"4abff6eb",
   918 => x"cff0c291",
   919 => x"e3c24abf",
   920 => x"a17248ea",
   921 => x"f2e3c278",
   922 => x"f978c048",
   923 => x"48c087e2",
   924 => x"e4e58ef4",
   925 => x"00000087",
   926 => x"ffffff00",
   927 => x"000e85ff",
   928 => x"000e8e00",
   929 => x"54414600",
   930 => x"20203233",
   931 => x"41460020",
   932 => x"20363154",
   933 => x"1e002020",
   934 => x"c348d4ff",
   935 => x"486878ff",
   936 => x"ff1e4f26",
   937 => x"ffc348d4",
   938 => x"48d0ff78",
   939 => x"ff78e1c8",
   940 => x"78d448d4",
   941 => x"48e7f0c2",
   942 => x"50bfd4ff",
   943 => x"ff1e4f26",
   944 => x"e0c048d0",
   945 => x"1e4f2678",
   946 => x"7087ccff",
   947 => x"c6029949",
   948 => x"a9fbc087",
   949 => x"7187f105",
   950 => x"0e4f2648",
   951 => x"0e5c5b5e",
   952 => x"4cc04b71",
   953 => x"7087f0fe",
   954 => x"c0029949",
   955 => x"ecc087f9",
   956 => x"f2c002a9",
   957 => x"a9fbc087",
   958 => x"87ebc002",
   959 => x"acb766cc",
   960 => x"d087c703",
   961 => x"87c20266",
   962 => x"99715371",
   963 => x"c187c202",
   964 => x"87c3fe84",
   965 => x"02994970",
   966 => x"ecc087cd",
   967 => x"87c702a9",
   968 => x"05a9fbc0",
   969 => x"d087d5ff",
   970 => x"87c30266",
   971 => x"c07b97c0",
   972 => x"c405a9ec",
   973 => x"c54a7487",
   974 => x"c04a7487",
   975 => x"48728a0a",
   976 => x"4d2687c2",
   977 => x"4b264c26",
   978 => x"fd1e4f26",
   979 => x"497087c9",
   980 => x"a9b7f0c0",
   981 => x"c087ca04",
   982 => x"01a9b7f9",
   983 => x"f0c087c3",
   984 => x"b7c1c189",
   985 => x"87ca04a9",
   986 => x"a9b7dac1",
   987 => x"c087c301",
   988 => x"487189f7",
   989 => x"5e0e4f26",
   990 => x"710e5c5b",
   991 => x"4cd4ff4a",
   992 => x"eac04972",
   993 => x"9b4b7087",
   994 => x"c187c202",
   995 => x"48d0ff8b",
   996 => x"c178c5c8",
   997 => x"49737cd5",
   998 => x"e2c231c6",
   999 => x"4abf97df",
  1000 => x"70b07148",
  1001 => x"48d0ff7c",
  1002 => x"487378c4",
  1003 => x"0e87d5fe",
  1004 => x"5d5c5b5e",
  1005 => x"7186f80e",
  1006 => x"fb7ec04c",
  1007 => x"4bc087e4",
  1008 => x"97dcc1c1",
  1009 => x"a9c049bf",
  1010 => x"fb87cf04",
  1011 => x"83c187f9",
  1012 => x"97dcc1c1",
  1013 => x"06ab49bf",
  1014 => x"c1c187f1",
  1015 => x"02bf97dc",
  1016 => x"f2fa87cf",
  1017 => x"99497087",
  1018 => x"c087c602",
  1019 => x"f105a9ec",
  1020 => x"fa4bc087",
  1021 => x"4d7087e1",
  1022 => x"c887dcfa",
  1023 => x"d6fa58a6",
  1024 => x"c14a7087",
  1025 => x"49a4c883",
  1026 => x"ad496997",
  1027 => x"c087c702",
  1028 => x"c005adff",
  1029 => x"a4c987e7",
  1030 => x"49699749",
  1031 => x"02a966c4",
  1032 => x"c04887c7",
  1033 => x"d405a8ff",
  1034 => x"49a4ca87",
  1035 => x"aa496997",
  1036 => x"c087c602",
  1037 => x"c405aaff",
  1038 => x"d07ec187",
  1039 => x"adecc087",
  1040 => x"c087c602",
  1041 => x"c405adfb",
  1042 => x"c14bc087",
  1043 => x"fe026e7e",
  1044 => x"e9f987e1",
  1045 => x"f8487387",
  1046 => x"87e6fb8e",
  1047 => x"5b5e0e00",
  1048 => x"1e0e5d5c",
  1049 => x"4cc04b71",
  1050 => x"c004ab4d",
  1051 => x"fec087e8",
  1052 => x"9d751eef",
  1053 => x"c087c402",
  1054 => x"c187c24a",
  1055 => x"f049724a",
  1056 => x"86c487df",
  1057 => x"84c17e70",
  1058 => x"87c2056e",
  1059 => x"85c14c73",
  1060 => x"ff06ac73",
  1061 => x"486e87d8",
  1062 => x"264d2626",
  1063 => x"264b264c",
  1064 => x"5b5e0e4f",
  1065 => x"1e0e5d5c",
  1066 => x"de494c71",
  1067 => x"c1f1c291",
  1068 => x"9785714d",
  1069 => x"ddc1026d",
  1070 => x"ecf0c287",
  1071 => x"82744abf",
  1072 => x"d8fe4972",
  1073 => x"6e7e7087",
  1074 => x"87f3c002",
  1075 => x"4bf4f0c2",
  1076 => x"49cb4a6e",
  1077 => x"87d0fffe",
  1078 => x"93cb4b74",
  1079 => x"83cae5c1",
  1080 => x"c4c183c4",
  1081 => x"49747bda",
  1082 => x"87c5c3c1",
  1083 => x"f1c27b75",
  1084 => x"49bf97c0",
  1085 => x"f4f0c21e",
  1086 => x"e4ddc149",
  1087 => x"7486c487",
  1088 => x"ecc2c149",
  1089 => x"c149c087",
  1090 => x"c287cbc4",
  1091 => x"c048e8f0",
  1092 => x"dd49c178",
  1093 => x"fd2687cb",
  1094 => x"6f4c87ff",
  1095 => x"6e696461",
  1096 => x"2e2e2e67",
  1097 => x"5b5e0e00",
  1098 => x"4b710e5c",
  1099 => x"ecf0c24a",
  1100 => x"497282bf",
  1101 => x"7087e6fc",
  1102 => x"c4029c4c",
  1103 => x"e8ec4987",
  1104 => x"ecf0c287",
  1105 => x"c178c048",
  1106 => x"87d5dc49",
  1107 => x"0e87ccfd",
  1108 => x"5d5c5b5e",
  1109 => x"c286f40e",
  1110 => x"c04df6e3",
  1111 => x"48a6c44c",
  1112 => x"f0c278c0",
  1113 => x"c049bfec",
  1114 => x"c1c106a9",
  1115 => x"f6e3c287",
  1116 => x"c0029848",
  1117 => x"fec087f8",
  1118 => x"66c81eef",
  1119 => x"c487c702",
  1120 => x"78c048a6",
  1121 => x"a6c487c5",
  1122 => x"c478c148",
  1123 => x"d0ec4966",
  1124 => x"7086c487",
  1125 => x"c484c14d",
  1126 => x"80c14866",
  1127 => x"c258a6c8",
  1128 => x"49bfecf0",
  1129 => x"87c603ac",
  1130 => x"ff059d75",
  1131 => x"4cc087c8",
  1132 => x"c3029d75",
  1133 => x"fec087e0",
  1134 => x"66c81eef",
  1135 => x"cc87c702",
  1136 => x"78c048a6",
  1137 => x"a6cc87c5",
  1138 => x"cc78c148",
  1139 => x"d0eb4966",
  1140 => x"7086c487",
  1141 => x"c2026e7e",
  1142 => x"496e87e9",
  1143 => x"699781cb",
  1144 => x"0299d049",
  1145 => x"c187d6c1",
  1146 => x"744ae5c4",
  1147 => x"c191cb49",
  1148 => x"7281cae5",
  1149 => x"c381c879",
  1150 => x"497451ff",
  1151 => x"f1c291de",
  1152 => x"85714dc1",
  1153 => x"7d97c1c2",
  1154 => x"c049a5c1",
  1155 => x"ecc251e0",
  1156 => x"02bf97c6",
  1157 => x"84c187d2",
  1158 => x"c24ba5c2",
  1159 => x"db4ac6ec",
  1160 => x"c3fafe49",
  1161 => x"87dbc187",
  1162 => x"c049a5cd",
  1163 => x"c284c151",
  1164 => x"4a6e4ba5",
  1165 => x"f9fe49cb",
  1166 => x"c6c187ee",
  1167 => x"e1c2c187",
  1168 => x"cb49744a",
  1169 => x"cae5c191",
  1170 => x"c2797281",
  1171 => x"bf97c6ec",
  1172 => x"7487d802",
  1173 => x"c191de49",
  1174 => x"c1f1c284",
  1175 => x"c283714b",
  1176 => x"dd4ac6ec",
  1177 => x"fff8fe49",
  1178 => x"7487d887",
  1179 => x"c293de4b",
  1180 => x"cb83c1f1",
  1181 => x"51c049a3",
  1182 => x"6e7384c1",
  1183 => x"fe49cb4a",
  1184 => x"c487e5f8",
  1185 => x"80c14866",
  1186 => x"c758a6c8",
  1187 => x"c5c003ac",
  1188 => x"fc056e87",
  1189 => x"487487e0",
  1190 => x"fcf78ef4",
  1191 => x"1e731e87",
  1192 => x"cb494b71",
  1193 => x"cae5c191",
  1194 => x"4aa1c881",
  1195 => x"48dfe2c2",
  1196 => x"a1c95012",
  1197 => x"dcc1c14a",
  1198 => x"ca501248",
  1199 => x"c0f1c281",
  1200 => x"c2501148",
  1201 => x"bf97c0f1",
  1202 => x"49c01e49",
  1203 => x"87d1d6c1",
  1204 => x"48e8f0c2",
  1205 => x"49c178de",
  1206 => x"2687c6d6",
  1207 => x"1e87fef6",
  1208 => x"cb494a71",
  1209 => x"cae5c191",
  1210 => x"1181c881",
  1211 => x"ecf0c248",
  1212 => x"ecf0c258",
  1213 => x"c178c048",
  1214 => x"87e5d549",
  1215 => x"c01e4f26",
  1216 => x"d1fcc049",
  1217 => x"1e4f2687",
  1218 => x"d2029971",
  1219 => x"dfe6c187",
  1220 => x"f750c048",
  1221 => x"dfcbc180",
  1222 => x"c3e5c140",
  1223 => x"c187ce78",
  1224 => x"c148dbe6",
  1225 => x"fc78fce4",
  1226 => x"fecbc180",
  1227 => x"0e4f2678",
  1228 => x"0e5c5b5e",
  1229 => x"cb4a4c71",
  1230 => x"cae5c192",
  1231 => x"49a2c882",
  1232 => x"974ba2c9",
  1233 => x"971e4b6b",
  1234 => x"ca1e4969",
  1235 => x"c0491282",
  1236 => x"c087cce7",
  1237 => x"87c9d449",
  1238 => x"f9c04974",
  1239 => x"8ef887d3",
  1240 => x"1e87f8f4",
  1241 => x"4b711e73",
  1242 => x"87c3ff49",
  1243 => x"fefe4973",
  1244 => x"87e9f487",
  1245 => x"711e731e",
  1246 => x"4aa3c64b",
  1247 => x"c187db02",
  1248 => x"87d6028a",
  1249 => x"dac1028a",
  1250 => x"c0028a87",
  1251 => x"028a87fc",
  1252 => x"8a87e1c0",
  1253 => x"c187cb02",
  1254 => x"49c787db",
  1255 => x"c187c0fd",
  1256 => x"f0c287de",
  1257 => x"c102bfec",
  1258 => x"c14887cb",
  1259 => x"f0f0c288",
  1260 => x"87c1c158",
  1261 => x"bff0f0c2",
  1262 => x"87f9c002",
  1263 => x"bfecf0c2",
  1264 => x"c280c148",
  1265 => x"c058f0f0",
  1266 => x"f0c287eb",
  1267 => x"c649bfec",
  1268 => x"f0f0c289",
  1269 => x"a9b7c059",
  1270 => x"c287da03",
  1271 => x"c048ecf0",
  1272 => x"c287d278",
  1273 => x"02bff0f0",
  1274 => x"f0c287cb",
  1275 => x"c648bfec",
  1276 => x"f0f0c280",
  1277 => x"d149c058",
  1278 => x"497387e7",
  1279 => x"87f1f6c0",
  1280 => x"0e87daf2",
  1281 => x"0e5c5b5e",
  1282 => x"66cc4c71",
  1283 => x"cb4b741e",
  1284 => x"cae5c193",
  1285 => x"4aa3c483",
  1286 => x"f2fe496a",
  1287 => x"cac187da",
  1288 => x"a3c87bdd",
  1289 => x"5166d449",
  1290 => x"d849a3c9",
  1291 => x"a3ca5166",
  1292 => x"5166dc49",
  1293 => x"87e3f126",
  1294 => x"5c5b5e0e",
  1295 => x"d0ff0e5d",
  1296 => x"59a6d886",
  1297 => x"c048a6c4",
  1298 => x"c180c478",
  1299 => x"c47866c4",
  1300 => x"c478c180",
  1301 => x"c278c180",
  1302 => x"c148f0f0",
  1303 => x"e8f0c278",
  1304 => x"a8de48bf",
  1305 => x"f387cb05",
  1306 => x"497087e5",
  1307 => x"ce59a6c8",
  1308 => x"ede887f8",
  1309 => x"87cfe987",
  1310 => x"7087dce8",
  1311 => x"acfbc04c",
  1312 => x"87d0c102",
  1313 => x"c10566d4",
  1314 => x"1ec087c2",
  1315 => x"c11ec11e",
  1316 => x"c01efde6",
  1317 => x"87ebfd49",
  1318 => x"4a66d0c1",
  1319 => x"496a82c4",
  1320 => x"517481c7",
  1321 => x"1ed81ec1",
  1322 => x"81c8496a",
  1323 => x"d887ece8",
  1324 => x"66c4c186",
  1325 => x"01a8c048",
  1326 => x"a6c487c7",
  1327 => x"ce78c148",
  1328 => x"66c4c187",
  1329 => x"cc88c148",
  1330 => x"87c358a6",
  1331 => x"cc87f8e7",
  1332 => x"78c248a6",
  1333 => x"cd029c74",
  1334 => x"66c487cc",
  1335 => x"66c8c148",
  1336 => x"c1cd03a8",
  1337 => x"48a6d887",
  1338 => x"eae678c0",
  1339 => x"c14c7087",
  1340 => x"c205acd0",
  1341 => x"66d887d6",
  1342 => x"87cee97e",
  1343 => x"a6dc4970",
  1344 => x"87d3e659",
  1345 => x"ecc04c70",
  1346 => x"eac105ac",
  1347 => x"4966c487",
  1348 => x"c0c191cb",
  1349 => x"a1c48166",
  1350 => x"c84d6a4a",
  1351 => x"66d84aa1",
  1352 => x"dfcbc152",
  1353 => x"87efe579",
  1354 => x"029c4c70",
  1355 => x"fbc087d8",
  1356 => x"87d202ac",
  1357 => x"dee55574",
  1358 => x"9c4c7087",
  1359 => x"c087c702",
  1360 => x"ff05acfb",
  1361 => x"e0c087ee",
  1362 => x"55c1c255",
  1363 => x"d47d97c0",
  1364 => x"a96e4966",
  1365 => x"c487db05",
  1366 => x"66c84866",
  1367 => x"87ca04a8",
  1368 => x"c14866c4",
  1369 => x"58a6c880",
  1370 => x"66c887c8",
  1371 => x"cc88c148",
  1372 => x"e2e458a6",
  1373 => x"c14c7087",
  1374 => x"c805acd0",
  1375 => x"4866d087",
  1376 => x"a6d480c1",
  1377 => x"acd0c158",
  1378 => x"87eafd02",
  1379 => x"d448a6dc",
  1380 => x"66d87866",
  1381 => x"a866dc48",
  1382 => x"87dcc905",
  1383 => x"48a6e0c0",
  1384 => x"c478f0c0",
  1385 => x"7866cc80",
  1386 => x"78c080c4",
  1387 => x"c048747e",
  1388 => x"f0c088fb",
  1389 => x"987058a6",
  1390 => x"87d7c802",
  1391 => x"c088cb48",
  1392 => x"7058a6f0",
  1393 => x"e9c00298",
  1394 => x"88c94887",
  1395 => x"58a6f0c0",
  1396 => x"c3029870",
  1397 => x"c44887e1",
  1398 => x"a6f0c088",
  1399 => x"02987058",
  1400 => x"c14887de",
  1401 => x"a6f0c088",
  1402 => x"02987058",
  1403 => x"c787c8c3",
  1404 => x"e0c087db",
  1405 => x"78c048a6",
  1406 => x"c14866cc",
  1407 => x"58a6d080",
  1408 => x"7087d4e2",
  1409 => x"acecc04c",
  1410 => x"c087d502",
  1411 => x"c60266e0",
  1412 => x"a6e4c087",
  1413 => x"7487c95c",
  1414 => x"88f0c048",
  1415 => x"58a6e8c0",
  1416 => x"02acecc0",
  1417 => x"eee187cc",
  1418 => x"c04c7087",
  1419 => x"ff05acec",
  1420 => x"e0c087f4",
  1421 => x"66d41e66",
  1422 => x"ecc01e49",
  1423 => x"e6c11e66",
  1424 => x"66d41efd",
  1425 => x"87fbf649",
  1426 => x"1eca1ec0",
  1427 => x"cb4966dc",
  1428 => x"66d8c191",
  1429 => x"48a6d881",
  1430 => x"d878a1c4",
  1431 => x"e149bf66",
  1432 => x"86d887f9",
  1433 => x"06a8b7c0",
  1434 => x"c187c7c1",
  1435 => x"c81ede1e",
  1436 => x"e149bf66",
  1437 => x"86c887e5",
  1438 => x"c0484970",
  1439 => x"e4c08808",
  1440 => x"b7c058a6",
  1441 => x"e9c006a8",
  1442 => x"66e0c087",
  1443 => x"a8b7dd48",
  1444 => x"6e87df03",
  1445 => x"e0c049bf",
  1446 => x"e0c08166",
  1447 => x"c1496651",
  1448 => x"81bf6e81",
  1449 => x"c051c1c2",
  1450 => x"c24966e0",
  1451 => x"81bf6e81",
  1452 => x"7ec151c0",
  1453 => x"e287dcc4",
  1454 => x"e4c087d0",
  1455 => x"c9e258a6",
  1456 => x"a6e8c087",
  1457 => x"a8ecc058",
  1458 => x"87cbc005",
  1459 => x"48a6e4c0",
  1460 => x"7866e0c0",
  1461 => x"ff87c4c0",
  1462 => x"c487fcde",
  1463 => x"91cb4966",
  1464 => x"4866c0c1",
  1465 => x"7e708071",
  1466 => x"82c84a6e",
  1467 => x"81ca496e",
  1468 => x"5166e0c0",
  1469 => x"4966e4c0",
  1470 => x"e0c081c1",
  1471 => x"48c18966",
  1472 => x"49703071",
  1473 => x"977189c1",
  1474 => x"ddf4c27a",
  1475 => x"e0c049bf",
  1476 => x"6a972966",
  1477 => x"9871484a",
  1478 => x"58a6f0c0",
  1479 => x"81c4496e",
  1480 => x"66dc4d69",
  1481 => x"a866d848",
  1482 => x"87c8c002",
  1483 => x"c048a6d8",
  1484 => x"87c5c078",
  1485 => x"c148a6d8",
  1486 => x"1e66d878",
  1487 => x"751ee0c0",
  1488 => x"d6deff49",
  1489 => x"7086c887",
  1490 => x"acb7c04c",
  1491 => x"87d4c106",
  1492 => x"e0c08574",
  1493 => x"75897449",
  1494 => x"dee1c14b",
  1495 => x"e5fe714a",
  1496 => x"85c287c6",
  1497 => x"4866e8c0",
  1498 => x"ecc080c1",
  1499 => x"ecc058a6",
  1500 => x"81c14966",
  1501 => x"c002a970",
  1502 => x"a6d887c8",
  1503 => x"c078c048",
  1504 => x"a6d887c5",
  1505 => x"d878c148",
  1506 => x"a4c21e66",
  1507 => x"48e0c049",
  1508 => x"49708871",
  1509 => x"ff49751e",
  1510 => x"c887c0dd",
  1511 => x"a8b7c086",
  1512 => x"87c0ff01",
  1513 => x"0266e8c0",
  1514 => x"6e87d1c0",
  1515 => x"c081c949",
  1516 => x"6e5166e8",
  1517 => x"efccc148",
  1518 => x"87ccc078",
  1519 => x"81c9496e",
  1520 => x"486e51c2",
  1521 => x"78e3cdc1",
  1522 => x"c6c07ec1",
  1523 => x"f6dbff87",
  1524 => x"6e4c7087",
  1525 => x"87f5c002",
  1526 => x"c84866c4",
  1527 => x"c004a866",
  1528 => x"66c487cb",
  1529 => x"c880c148",
  1530 => x"e0c058a6",
  1531 => x"4866c887",
  1532 => x"a6cc88c1",
  1533 => x"87d5c058",
  1534 => x"05acc6c1",
  1535 => x"cc87c8c0",
  1536 => x"80c14866",
  1537 => x"ff58a6d0",
  1538 => x"7087fcda",
  1539 => x"4866d04c",
  1540 => x"a6d480c1",
  1541 => x"029c7458",
  1542 => x"c487cbc0",
  1543 => x"c8c14866",
  1544 => x"f204a866",
  1545 => x"daff87ff",
  1546 => x"66c487d4",
  1547 => x"03a8c748",
  1548 => x"c287e5c0",
  1549 => x"c048f0f0",
  1550 => x"4966c478",
  1551 => x"c0c191cb",
  1552 => x"a1c48166",
  1553 => x"c04a6a4a",
  1554 => x"66c47952",
  1555 => x"c880c148",
  1556 => x"a8c758a6",
  1557 => x"87dbff04",
  1558 => x"e08ed0ff",
  1559 => x"203a87fb",
  1560 => x"1e731e00",
  1561 => x"029b4b71",
  1562 => x"f0c287c6",
  1563 => x"78c048ec",
  1564 => x"f0c21ec7",
  1565 => x"1e49bfec",
  1566 => x"1ecae5c1",
  1567 => x"bfe8f0c2",
  1568 => x"87f4ee49",
  1569 => x"f0c286cc",
  1570 => x"e949bfe8",
  1571 => x"9b7387f9",
  1572 => x"c187c802",
  1573 => x"c049cae5",
  1574 => x"ff87e8e5",
  1575 => x"1e87fedf",
  1576 => x"48dfe2c2",
  1577 => x"e6c150c0",
  1578 => x"c049bfed",
  1579 => x"c087c5fb",
  1580 => x"1e4f2648",
  1581 => x"c187e5c7",
  1582 => x"87e5fe49",
  1583 => x"87e0e9fe",
  1584 => x"cd029870",
  1585 => x"ddf2fe87",
  1586 => x"02987087",
  1587 => x"4ac187c4",
  1588 => x"4ac087c2",
  1589 => x"ce059a72",
  1590 => x"c11ec087",
  1591 => x"c049c3e4",
  1592 => x"c487eff0",
  1593 => x"c087fe86",
  1594 => x"cee4c11e",
  1595 => x"e1f0c049",
  1596 => x"fe1ec087",
  1597 => x"497087e9",
  1598 => x"87d6f0c0",
  1599 => x"f887dcc3",
  1600 => x"534f268e",
  1601 => x"61662044",
  1602 => x"64656c69",
  1603 => x"6f42002e",
  1604 => x"6e69746f",
  1605 => x"2e2e2e67",
  1606 => x"e8c01e00",
  1607 => x"f3c087c1",
  1608 => x"87f687e6",
  1609 => x"c21e4f26",
  1610 => x"c048ecf0",
  1611 => x"e8f0c278",
  1612 => x"fd78c048",
  1613 => x"87e187fd",
  1614 => x"4f2648c0",
  1615 => x"78452080",
  1616 => x"80007469",
  1617 => x"63614220",
  1618 => x"12df006b",
  1619 => x"2c410000",
  1620 => x"00000000",
  1621 => x"0012df00",
  1622 => x"002c5f00",
  1623 => x"00000000",
  1624 => x"000012df",
  1625 => x"00002c7d",
  1626 => x"df000000",
  1627 => x"9b000012",
  1628 => x"0000002c",
  1629 => x"12df0000",
  1630 => x"2cb90000",
  1631 => x"00000000",
  1632 => x"0012df00",
  1633 => x"002cd700",
  1634 => x"00000000",
  1635 => x"000012df",
  1636 => x"00002cf5",
  1637 => x"df000000",
  1638 => x"00000012",
  1639 => x"00000000",
  1640 => x"13740000",
  1641 => x"00000000",
  1642 => x"00000000",
  1643 => x"0019b100",
  1644 => x"4f4f4200",
  1645 => x"20202054",
  1646 => x"4d4f5220",
  1647 => x"616f4c00",
  1648 => x"2e2a2064",
  1649 => x"f0fe1e00",
  1650 => x"cd78c048",
  1651 => x"26097909",
  1652 => x"fe1e1e4f",
  1653 => x"487ebff0",
  1654 => x"1e4f2626",
  1655 => x"c148f0fe",
  1656 => x"1e4f2678",
  1657 => x"c048f0fe",
  1658 => x"1e4f2678",
  1659 => x"52c04a71",
  1660 => x"0e4f2652",
  1661 => x"5d5c5b5e",
  1662 => x"7186f40e",
  1663 => x"7e6d974d",
  1664 => x"974ca5c1",
  1665 => x"a6c8486c",
  1666 => x"c4486e58",
  1667 => x"c505a866",
  1668 => x"c048ff87",
  1669 => x"caff87e6",
  1670 => x"49a5c287",
  1671 => x"714b6c97",
  1672 => x"6b974ba3",
  1673 => x"7e6c974b",
  1674 => x"80c1486e",
  1675 => x"c758a6c8",
  1676 => x"58a6cc98",
  1677 => x"fe7c9770",
  1678 => x"487387e1",
  1679 => x"4d268ef4",
  1680 => x"4b264c26",
  1681 => x"5e0e4f26",
  1682 => x"f40e5c5b",
  1683 => x"d84c7186",
  1684 => x"ffc34a66",
  1685 => x"4ba4c29a",
  1686 => x"73496c97",
  1687 => x"517249a1",
  1688 => x"6e7e6c97",
  1689 => x"c880c148",
  1690 => x"98c758a6",
  1691 => x"7058a6cc",
  1692 => x"ff8ef454",
  1693 => x"1e1e87ca",
  1694 => x"e087e8fd",
  1695 => x"c0494abf",
  1696 => x"0299c0e0",
  1697 => x"1e7287cb",
  1698 => x"49d3f4c2",
  1699 => x"c487f7fe",
  1700 => x"87fdfc86",
  1701 => x"c2fd7e70",
  1702 => x"4f262687",
  1703 => x"d3f4c21e",
  1704 => x"87c7fd49",
  1705 => x"49f6e9c1",
  1706 => x"c587dafc",
  1707 => x"4f2687d9",
  1708 => x"5c5b5e0e",
  1709 => x"f4c20e5d",
  1710 => x"c14abff2",
  1711 => x"49bfc4ec",
  1712 => x"71bc724c",
  1713 => x"87dbfc4d",
  1714 => x"49744bc0",
  1715 => x"d50299d0",
  1716 => x"d0497587",
  1717 => x"c01e7199",
  1718 => x"d6f2c11e",
  1719 => x"1282734a",
  1720 => x"87e4c049",
  1721 => x"2cc186c8",
  1722 => x"abc8832d",
  1723 => x"87daff04",
  1724 => x"c187e8fb",
  1725 => x"c248c4ec",
  1726 => x"78bff2f4",
  1727 => x"4c264d26",
  1728 => x"4f264b26",
  1729 => x"00000000",
  1730 => x"48d0ff1e",
  1731 => x"ff78e1c8",
  1732 => x"78c548d4",
  1733 => x"c30266c4",
  1734 => x"78e0c387",
  1735 => x"c60266c8",
  1736 => x"48d4ff87",
  1737 => x"ff78f0c3",
  1738 => x"787148d4",
  1739 => x"c848d0ff",
  1740 => x"e0c078e1",
  1741 => x"0e4f2678",
  1742 => x"0e5c5b5e",
  1743 => x"f4c24c71",
  1744 => x"eefa49d3",
  1745 => x"c04a7087",
  1746 => x"c204aab7",
  1747 => x"e0c387e3",
  1748 => x"87c905aa",
  1749 => x"48faefc1",
  1750 => x"d4c278c1",
  1751 => x"aaf0c387",
  1752 => x"c187c905",
  1753 => x"c148f6ef",
  1754 => x"87f5c178",
  1755 => x"bffaefc1",
  1756 => x"7287c702",
  1757 => x"b3c0c24b",
  1758 => x"4b7287c2",
  1759 => x"d1059c74",
  1760 => x"f6efc187",
  1761 => x"efc11ebf",
  1762 => x"721ebffa",
  1763 => x"87f8fd49",
  1764 => x"efc186c8",
  1765 => x"c002bff6",
  1766 => x"497387e0",
  1767 => x"9129b7c4",
  1768 => x"81d6f1c1",
  1769 => x"9acf4a73",
  1770 => x"48c192c2",
  1771 => x"4a703072",
  1772 => x"4872baff",
  1773 => x"79709869",
  1774 => x"497387db",
  1775 => x"9129b7c4",
  1776 => x"81d6f1c1",
  1777 => x"9acf4a73",
  1778 => x"48c392c2",
  1779 => x"4a703072",
  1780 => x"70b06948",
  1781 => x"faefc179",
  1782 => x"c178c048",
  1783 => x"c048f6ef",
  1784 => x"d3f4c278",
  1785 => x"87cbf849",
  1786 => x"b7c04a70",
  1787 => x"ddfd03aa",
  1788 => x"fc48c087",
  1789 => x"000087c8",
  1790 => x"00000000",
  1791 => x"711e0000",
  1792 => x"f2fc494a",
  1793 => x"1e4f2687",
  1794 => x"49724ac0",
  1795 => x"f1c191c4",
  1796 => x"79c081d6",
  1797 => x"b7d082c1",
  1798 => x"87ee04aa",
  1799 => x"5e0e4f26",
  1800 => x"0e5d5c5b",
  1801 => x"faf64d71",
  1802 => x"c44a7587",
  1803 => x"c1922ab7",
  1804 => x"7582d6f1",
  1805 => x"c29ccf4c",
  1806 => x"4b496a94",
  1807 => x"9bc32b74",
  1808 => x"307448c2",
  1809 => x"bcff4c70",
  1810 => x"98714874",
  1811 => x"caf67a70",
  1812 => x"fa487387",
  1813 => x"000087e6",
  1814 => x"00000000",
  1815 => x"00000000",
  1816 => x"00000000",
  1817 => x"00000000",
  1818 => x"00000000",
  1819 => x"00000000",
  1820 => x"00000000",
  1821 => x"00000000",
  1822 => x"00000000",
  1823 => x"00000000",
  1824 => x"00000000",
  1825 => x"00000000",
  1826 => x"00000000",
  1827 => x"00000000",
  1828 => x"00000000",
  1829 => x"1e160000",
  1830 => x"362e2526",
  1831 => x"ff1e3e3d",
  1832 => x"e1c848d0",
  1833 => x"ff487178",
  1834 => x"267808d4",
  1835 => x"d0ff1e4f",
  1836 => x"78e1c848",
  1837 => x"d4ff4871",
  1838 => x"66c47808",
  1839 => x"08d4ff48",
  1840 => x"1e4f2678",
  1841 => x"66c44a71",
  1842 => x"49721e49",
  1843 => x"ff87deff",
  1844 => x"e0c048d0",
  1845 => x"4f262678",
  1846 => x"c24a711e",
  1847 => x"c303aab7",
  1848 => x"87c28287",
  1849 => x"66c482ce",
  1850 => x"ff49721e",
  1851 => x"262687d5",
  1852 => x"d4ff1e4f",
  1853 => x"7affc34a",
  1854 => x"c848d0ff",
  1855 => x"7ade78e1",
  1856 => x"bfddf4c2",
  1857 => x"c848497a",
  1858 => x"717a7028",
  1859 => x"7028d048",
  1860 => x"d848717a",
  1861 => x"ff7a7028",
  1862 => x"e0c048d0",
  1863 => x"0e4f2678",
  1864 => x"5d5c5b5e",
  1865 => x"c24c710e",
  1866 => x"4dbfddf4",
  1867 => x"d02b744b",
  1868 => x"83c19b66",
  1869 => x"04ab66d4",
  1870 => x"4bc087c2",
  1871 => x"66d04a74",
  1872 => x"ff317249",
  1873 => x"739975b9",
  1874 => x"70307248",
  1875 => x"b071484a",
  1876 => x"58e1f4c2",
  1877 => x"2687dafe",
  1878 => x"264c264d",
  1879 => x"1e4f264b",
  1880 => x"c848d0ff",
  1881 => x"487178c9",
  1882 => x"7808d4ff",
  1883 => x"711e4f26",
  1884 => x"87eb494a",
  1885 => x"c848d0ff",
  1886 => x"1e4f2678",
  1887 => x"4b711e73",
  1888 => x"bfedf4c2",
  1889 => x"c287c302",
  1890 => x"d0ff87eb",
  1891 => x"78c9c848",
  1892 => x"e0c04973",
  1893 => x"48d4ffb1",
  1894 => x"f4c27871",
  1895 => x"78c048e1",
  1896 => x"c50266c8",
  1897 => x"49ffc387",
  1898 => x"49c087c2",
  1899 => x"59e9f4c2",
  1900 => x"c60266cc",
  1901 => x"d5d5c587",
  1902 => x"cf87c44a",
  1903 => x"c24affff",
  1904 => x"c25aedf4",
  1905 => x"c148edf4",
  1906 => x"2687c478",
  1907 => x"264c264d",
  1908 => x"0e4f264b",
  1909 => x"5d5c5b5e",
  1910 => x"c24a710e",
  1911 => x"4cbfe9f4",
  1912 => x"cb029a72",
  1913 => x"91c84987",
  1914 => x"4bf1f5c1",
  1915 => x"87c48371",
  1916 => x"4bf1f9c1",
  1917 => x"49134dc0",
  1918 => x"f4c29974",
  1919 => x"ffb9bfe5",
  1920 => x"787148d4",
  1921 => x"852cb7c1",
  1922 => x"04adb7c8",
  1923 => x"f4c287e8",
  1924 => x"c848bfe1",
  1925 => x"e5f4c280",
  1926 => x"87effe58",
  1927 => x"711e731e",
  1928 => x"9a4a134b",
  1929 => x"7287cb02",
  1930 => x"87e7fe49",
  1931 => x"059a4a13",
  1932 => x"dafe87f5",
  1933 => x"f4c21e87",
  1934 => x"c249bfe1",
  1935 => x"c148e1f4",
  1936 => x"c0c478a1",
  1937 => x"db03a9b7",
  1938 => x"48d4ff87",
  1939 => x"bfe5f4c2",
  1940 => x"e1f4c278",
  1941 => x"f4c249bf",
  1942 => x"a1c148e1",
  1943 => x"b7c0c478",
  1944 => x"87e504a9",
  1945 => x"c848d0ff",
  1946 => x"edf4c278",
  1947 => x"2678c048",
  1948 => x"0000004f",
  1949 => x"00000000",
  1950 => x"00000000",
  1951 => x"00005f5f",
  1952 => x"03030000",
  1953 => x"00030300",
  1954 => x"7f7f1400",
  1955 => x"147f7f14",
  1956 => x"2e240000",
  1957 => x"123a6b6b",
  1958 => x"366a4c00",
  1959 => x"32566c18",
  1960 => x"4f7e3000",
  1961 => x"683a7759",
  1962 => x"04000040",
  1963 => x"00000307",
  1964 => x"1c000000",
  1965 => x"0041633e",
  1966 => x"41000000",
  1967 => x"001c3e63",
  1968 => x"3e2a0800",
  1969 => x"2a3e1c1c",
  1970 => x"08080008",
  1971 => x"08083e3e",
  1972 => x"80000000",
  1973 => x"000060e0",
  1974 => x"08080000",
  1975 => x"08080808",
  1976 => x"00000000",
  1977 => x"00006060",
  1978 => x"30604000",
  1979 => x"03060c18",
  1980 => x"7f3e0001",
  1981 => x"3e7f4d59",
  1982 => x"06040000",
  1983 => x"00007f7f",
  1984 => x"63420000",
  1985 => x"464f5971",
  1986 => x"63220000",
  1987 => x"367f4949",
  1988 => x"161c1800",
  1989 => x"107f7f13",
  1990 => x"67270000",
  1991 => x"397d4545",
  1992 => x"7e3c0000",
  1993 => x"3079494b",
  1994 => x"01010000",
  1995 => x"070f7971",
  1996 => x"7f360000",
  1997 => x"367f4949",
  1998 => x"4f060000",
  1999 => x"1e3f6949",
  2000 => x"00000000",
  2001 => x"00006666",
  2002 => x"80000000",
  2003 => x"000066e6",
  2004 => x"08080000",
  2005 => x"22221414",
  2006 => x"14140000",
  2007 => x"14141414",
  2008 => x"22220000",
  2009 => x"08081414",
  2010 => x"03020000",
  2011 => x"060f5951",
  2012 => x"417f3e00",
  2013 => x"1e1f555d",
  2014 => x"7f7e0000",
  2015 => x"7e7f0909",
  2016 => x"7f7f0000",
  2017 => x"367f4949",
  2018 => x"3e1c0000",
  2019 => x"41414163",
  2020 => x"7f7f0000",
  2021 => x"1c3e6341",
  2022 => x"7f7f0000",
  2023 => x"41414949",
  2024 => x"7f7f0000",
  2025 => x"01010909",
  2026 => x"7f3e0000",
  2027 => x"7a7b4941",
  2028 => x"7f7f0000",
  2029 => x"7f7f0808",
  2030 => x"41000000",
  2031 => x"00417f7f",
  2032 => x"60200000",
  2033 => x"3f7f4040",
  2034 => x"087f7f00",
  2035 => x"4163361c",
  2036 => x"7f7f0000",
  2037 => x"40404040",
  2038 => x"067f7f00",
  2039 => x"7f7f060c",
  2040 => x"067f7f00",
  2041 => x"7f7f180c",
  2042 => x"7f3e0000",
  2043 => x"3e7f4141",
  2044 => x"7f7f0000",
  2045 => x"060f0909",
  2046 => x"417f3e00",
  2047 => x"407e7f61",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
