library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"7f7f0000",
     1 => x"667f1909",
     2 => x"6f260000",
     3 => x"327b594d",
     4 => x"01010000",
     5 => x"01017f7f",
     6 => x"7f3f0000",
     7 => x"3f7f4040",
     8 => x"3f0f0000",
     9 => x"0f3f7070",
    10 => x"307f7f00",
    11 => x"7f7f3018",
    12 => x"36634100",
    13 => x"63361c1c",
    14 => x"06030141",
    15 => x"03067c7c",
    16 => x"59716101",
    17 => x"4143474d",
    18 => x"7f000000",
    19 => x"0041417f",
    20 => x"06030100",
    21 => x"6030180c",
    22 => x"41000040",
    23 => x"007f7f41",
    24 => x"060c0800",
    25 => x"080c0603",
    26 => x"80808000",
    27 => x"80808080",
    28 => x"00000000",
    29 => x"00040703",
    30 => x"74200000",
    31 => x"787c5454",
    32 => x"7f7f0000",
    33 => x"387c4444",
    34 => x"7c380000",
    35 => x"00444444",
    36 => x"7c380000",
    37 => x"7f7f4444",
    38 => x"7c380000",
    39 => x"185c5454",
    40 => x"7e040000",
    41 => x"0005057f",
    42 => x"bc180000",
    43 => x"7cfca4a4",
    44 => x"7f7f0000",
    45 => x"787c0404",
    46 => x"00000000",
    47 => x"00407d3d",
    48 => x"80800000",
    49 => x"007dfd80",
    50 => x"7f7f0000",
    51 => x"446c3810",
    52 => x"00000000",
    53 => x"00407f3f",
    54 => x"0c7c7c00",
    55 => x"787c0c18",
    56 => x"7c7c0000",
    57 => x"787c0404",
    58 => x"7c380000",
    59 => x"387c4444",
    60 => x"fcfc0000",
    61 => x"183c2424",
    62 => x"3c180000",
    63 => x"fcfc2424",
    64 => x"7c7c0000",
    65 => x"080c0404",
    66 => x"5c480000",
    67 => x"20745454",
    68 => x"3f040000",
    69 => x"0044447f",
    70 => x"7c3c0000",
    71 => x"7c7c4040",
    72 => x"3c1c0000",
    73 => x"1c3c6060",
    74 => x"607c3c00",
    75 => x"3c7c6030",
    76 => x"386c4400",
    77 => x"446c3810",
    78 => x"bc1c0000",
    79 => x"1c3c60e0",
    80 => x"64440000",
    81 => x"444c5c74",
    82 => x"08080000",
    83 => x"4141773e",
    84 => x"00000000",
    85 => x"00007f7f",
    86 => x"41410000",
    87 => x"08083e77",
    88 => x"01010200",
    89 => x"01020203",
    90 => x"7f7f7f00",
    91 => x"7f7f7f7f",
    92 => x"1c080800",
    93 => x"7f3e3e1c",
    94 => x"3e7f7f7f",
    95 => x"081c1c3e",
    96 => x"18100008",
    97 => x"10187c7c",
    98 => x"30100000",
    99 => x"10307c7c",
   100 => x"60301000",
   101 => x"061e7860",
   102 => x"3c664200",
   103 => x"42663c18",
   104 => x"6a387800",
   105 => x"386cc6c2",
   106 => x"00006000",
   107 => x"60000060",
   108 => x"5b5e0e00",
   109 => x"1e0e5d5c",
   110 => x"f4c24c71",
   111 => x"c04dbffe",
   112 => x"741ec04b",
   113 => x"87c702ab",
   114 => x"c048a6c4",
   115 => x"c487c578",
   116 => x"78c148a6",
   117 => x"731e66c4",
   118 => x"87dfee49",
   119 => x"e0c086c8",
   120 => x"87efef49",
   121 => x"6a4aa5c4",
   122 => x"87f0f049",
   123 => x"cb87c6f1",
   124 => x"c883c185",
   125 => x"ff04abb7",
   126 => x"262687c7",
   127 => x"264c264d",
   128 => x"1e4f264b",
   129 => x"f5c24a71",
   130 => x"f5c25ac2",
   131 => x"78c748c2",
   132 => x"87ddfe49",
   133 => x"731e4f26",
   134 => x"c04a711e",
   135 => x"d303aab7",
   136 => x"e7d5c287",
   137 => x"87c405bf",
   138 => x"87c24bc1",
   139 => x"d5c24bc0",
   140 => x"87c45beb",
   141 => x"5aebd5c2",
   142 => x"bfe7d5c2",
   143 => x"c19ac14a",
   144 => x"ec49a2c0",
   145 => x"48fc87e8",
   146 => x"bfe7d5c2",
   147 => x"87effe78",
   148 => x"c44a711e",
   149 => x"49721e66",
   150 => x"2687fde9",
   151 => x"c21e4f26",
   152 => x"49bfe7d5",
   153 => x"c287d7e6",
   154 => x"e848f6f4",
   155 => x"f4c278bf",
   156 => x"bfec48f2",
   157 => x"f6f4c278",
   158 => x"c3494abf",
   159 => x"b7c899ff",
   160 => x"7148722a",
   161 => x"fef4c2b0",
   162 => x"0e4f2658",
   163 => x"5d5c5b5e",
   164 => x"ff4b710e",
   165 => x"f4c287c8",
   166 => x"50c048f1",
   167 => x"fde54973",
   168 => x"4c497087",
   169 => x"eecb9cc2",
   170 => x"87c3cb49",
   171 => x"c24d4970",
   172 => x"bf97f1f4",
   173 => x"87e2c105",
   174 => x"c24966d0",
   175 => x"99bffaf4",
   176 => x"d487d605",
   177 => x"f4c24966",
   178 => x"0599bff2",
   179 => x"497387cb",
   180 => x"7087cbe5",
   181 => x"c1c10298",
   182 => x"fe4cc187",
   183 => x"497587c0",
   184 => x"7087d8ca",
   185 => x"87c60298",
   186 => x"48f1f4c2",
   187 => x"f4c250c1",
   188 => x"05bf97f1",
   189 => x"c287e3c0",
   190 => x"49bffaf4",
   191 => x"059966d0",
   192 => x"c287d6ff",
   193 => x"49bff2f4",
   194 => x"059966d4",
   195 => x"7387caff",
   196 => x"87cae449",
   197 => x"fe059870",
   198 => x"487487ff",
   199 => x"0e87dcfb",
   200 => x"5d5c5b5e",
   201 => x"c086f40e",
   202 => x"bfec4c4d",
   203 => x"48a6c47e",
   204 => x"bffef4c2",
   205 => x"c01ec178",
   206 => x"fd49c71e",
   207 => x"86c887cd",
   208 => x"cd029870",
   209 => x"fb49ff87",
   210 => x"dac187cc",
   211 => x"87cee349",
   212 => x"f4c24dc1",
   213 => x"02bf97f1",
   214 => x"c3d587c3",
   215 => x"f6f4c287",
   216 => x"d5c24bbf",
   217 => x"c005bfe7",
   218 => x"fdc387e9",
   219 => x"87eee249",
   220 => x"e249fac3",
   221 => x"497387e8",
   222 => x"7199ffc3",
   223 => x"fb49c01e",
   224 => x"497387ce",
   225 => x"7129b7c8",
   226 => x"fb49c11e",
   227 => x"86c887c2",
   228 => x"c287fac5",
   229 => x"4bbffaf4",
   230 => x"87dd029b",
   231 => x"bfe3d5c2",
   232 => x"87d7c749",
   233 => x"c4059870",
   234 => x"d24bc087",
   235 => x"49e0c287",
   236 => x"c287fcc6",
   237 => x"c658e7d5",
   238 => x"e3d5c287",
   239 => x"7378c048",
   240 => x"0599c249",
   241 => x"ebc387cd",
   242 => x"87d2e149",
   243 => x"99c24970",
   244 => x"fb87c202",
   245 => x"c149734c",
   246 => x"87cd0599",
   247 => x"e049f4c3",
   248 => x"497087fc",
   249 => x"c20299c2",
   250 => x"734cfa87",
   251 => x"0599c849",
   252 => x"f5c387cd",
   253 => x"87e6e049",
   254 => x"99c24970",
   255 => x"c287d402",
   256 => x"02bfc2f5",
   257 => x"c14887c9",
   258 => x"c6f5c288",
   259 => x"ff87c258",
   260 => x"734dc14c",
   261 => x"0599c449",
   262 => x"f2c387ce",
   263 => x"fddfff49",
   264 => x"c2497087",
   265 => x"87db0299",
   266 => x"bfc2f5c2",
   267 => x"b7c7487e",
   268 => x"87cb03a8",
   269 => x"80c1486e",
   270 => x"58c6f5c2",
   271 => x"fe87c2c0",
   272 => x"c34dc14c",
   273 => x"dfff49fd",
   274 => x"497087d4",
   275 => x"d50299c2",
   276 => x"c2f5c287",
   277 => x"c9c002bf",
   278 => x"c2f5c287",
   279 => x"c078c048",
   280 => x"4cfd87c2",
   281 => x"fac34dc1",
   282 => x"f1deff49",
   283 => x"c2497087",
   284 => x"87d90299",
   285 => x"bfc2f5c2",
   286 => x"a8b7c748",
   287 => x"87c9c003",
   288 => x"48c2f5c2",
   289 => x"c2c078c7",
   290 => x"c14cfc87",
   291 => x"acb7c04d",
   292 => x"87d1c003",
   293 => x"c14a66c4",
   294 => x"026a82d8",
   295 => x"6a87c6c0",
   296 => x"7349744b",
   297 => x"c31ec00f",
   298 => x"dac11ef0",
   299 => x"87dbf749",
   300 => x"987086c8",
   301 => x"87e2c002",
   302 => x"c248a6c8",
   303 => x"78bfc2f5",
   304 => x"cb4966c8",
   305 => x"4866c491",
   306 => x"7e708071",
   307 => x"c002bf6e",
   308 => x"bf6e87c8",
   309 => x"4966c84b",
   310 => x"9d750f73",
   311 => x"87c8c002",
   312 => x"bfc2f5c2",
   313 => x"87c9f349",
   314 => x"bfebd5c2",
   315 => x"87ddc002",
   316 => x"87c7c249",
   317 => x"c0029870",
   318 => x"f5c287d3",
   319 => x"f249bfc2",
   320 => x"49c087ef",
   321 => x"c287cff4",
   322 => x"c048ebd5",
   323 => x"f38ef478",
   324 => x"5e0e87e9",
   325 => x"0e5d5c5b",
   326 => x"c24c711e",
   327 => x"49bffef4",
   328 => x"4da1cdc1",
   329 => x"6981d1c1",
   330 => x"029c747e",
   331 => x"a5c487cf",
   332 => x"c27b744b",
   333 => x"49bffef4",
   334 => x"6e87c8f3",
   335 => x"059c747b",
   336 => x"4bc087c4",
   337 => x"4bc187c2",
   338 => x"c9f34973",
   339 => x"0266d487",
   340 => x"da4987c7",
   341 => x"c24a7087",
   342 => x"c24ac087",
   343 => x"265aefd5",
   344 => x"0087d8f2",
   345 => x"00000000",
   346 => x"00000000",
   347 => x"1e000000",
   348 => x"c8ff4a71",
   349 => x"a17249bf",
   350 => x"1e4f2648",
   351 => x"89bfc8ff",
   352 => x"c0c0c0fe",
   353 => x"01a9c0c0",
   354 => x"4ac087c4",
   355 => x"4ac187c2",
   356 => x"4f264872",
   357 => x"5c5b5e0e",
   358 => x"4b710e5d",
   359 => x"d04cd4ff",
   360 => x"78c04866",
   361 => x"dbff49d6",
   362 => x"ffc387f4",
   363 => x"c3496c7c",
   364 => x"4d7199ff",
   365 => x"99f0c349",
   366 => x"05a9e0c1",
   367 => x"ffc387cb",
   368 => x"c3486c7c",
   369 => x"0866d098",
   370 => x"7cffc378",
   371 => x"c8494a6c",
   372 => x"7cffc331",
   373 => x"b2714a6c",
   374 => x"31c84972",
   375 => x"6c7cffc3",
   376 => x"72b2714a",
   377 => x"c331c849",
   378 => x"4a6c7cff",
   379 => x"d0ffb271",
   380 => x"78e0c048",
   381 => x"c2029b73",
   382 => x"757b7287",
   383 => x"264d2648",
   384 => x"264b264c",
   385 => x"4f261e4f",
   386 => x"5c5b5e0e",
   387 => x"7686f80e",
   388 => x"49a6c81e",
   389 => x"c487fdfd",
   390 => x"6e4b7086",
   391 => x"03a8c448",
   392 => x"7387cac3",
   393 => x"9af0c34a",
   394 => x"02aad0c1",
   395 => x"e0c187c7",
   396 => x"f8c205aa",
   397 => x"c8497387",
   398 => x"87c30299",
   399 => x"7387c6ff",
   400 => x"c29cc34c",
   401 => x"cfc105ac",
   402 => x"4966c487",
   403 => x"1e7131c9",
   404 => x"c14a66c4",
   405 => x"f5c292c8",
   406 => x"817249c6",
   407 => x"87efd2fe",
   408 => x"1e4966c4",
   409 => x"ff49e3c0",
   410 => x"d887d8d9",
   411 => x"edd8ff49",
   412 => x"1ec0c887",
   413 => x"49f6e3c2",
   414 => x"87c4ebfd",
   415 => x"c048d0ff",
   416 => x"e3c278e0",
   417 => x"66d01ef6",
   418 => x"92c8c14a",
   419 => x"49c6f5c2",
   420 => x"cdfe8172",
   421 => x"86d087f7",
   422 => x"c105acc1",
   423 => x"66c487cf",
   424 => x"7131c949",
   425 => x"4a66c41e",
   426 => x"c292c8c1",
   427 => x"7249c6f5",
   428 => x"dad1fe81",
   429 => x"f6e3c287",
   430 => x"4a66c81e",
   431 => x"c292c8c1",
   432 => x"7249c6f5",
   433 => x"c1ccfe81",
   434 => x"4966c887",
   435 => x"49e3c01e",
   436 => x"87efd7ff",
   437 => x"d7ff49d7",
   438 => x"c0c887c4",
   439 => x"f6e3c21e",
   440 => x"c5e9fd49",
   441 => x"ff86d087",
   442 => x"e0c048d0",
   443 => x"fc8ef878",
   444 => x"5e0e87cd",
   445 => x"0e5d5c5b",
   446 => x"ff4d711e",
   447 => x"66d44cd4",
   448 => x"b7c3487e",
   449 => x"87c506a8",
   450 => x"e3c148c0",
   451 => x"fe497587",
   452 => x"7587e3e1",
   453 => x"4b66c41e",
   454 => x"c293c8c1",
   455 => x"7383c6f5",
   456 => x"cfc6fe49",
   457 => x"6b83c887",
   458 => x"48d0ff4b",
   459 => x"dd78e1c8",
   460 => x"c349737c",
   461 => x"7c7199ff",
   462 => x"b7c84973",
   463 => x"99ffc329",
   464 => x"49737c71",
   465 => x"c329b7d0",
   466 => x"7c7199ff",
   467 => x"b7d84973",
   468 => x"c07c7129",
   469 => x"7c7c7c7c",
   470 => x"7c7c7c7c",
   471 => x"7c7c7c7c",
   472 => x"c478e0c0",
   473 => x"49dc1e66",
   474 => x"87d7d5ff",
   475 => x"487386c8",
   476 => x"87c9fa26",
   477 => x"5c5b5e0e",
   478 => x"711e0e5d",
   479 => x"4bd4ff7e",
   480 => x"f9c21e6e",
   481 => x"c4fe49e6",
   482 => x"86c487ea",
   483 => x"029d4d70",
   484 => x"c287c3c3",
   485 => x"4cbfeef9",
   486 => x"dffe496e",
   487 => x"d0ff87d8",
   488 => x"78c5c848",
   489 => x"c07bd6c1",
   490 => x"c17b154a",
   491 => x"b7e0c082",
   492 => x"87f504aa",
   493 => x"c448d0ff",
   494 => x"78c5c878",
   495 => x"c17bd3c1",
   496 => x"7478c47b",
   497 => x"fcc1029c",
   498 => x"f6e3c287",
   499 => x"4dc0c87e",
   500 => x"acb7c08c",
   501 => x"c887c603",
   502 => x"c04da4c0",
   503 => x"e7f0c24c",
   504 => x"d049bf97",
   505 => x"87d20299",
   506 => x"f9c21ec0",
   507 => x"c7fe49e6",
   508 => x"86c487d8",
   509 => x"c04a4970",
   510 => x"e3c287ef",
   511 => x"f9c21ef6",
   512 => x"c7fe49e6",
   513 => x"86c487c4",
   514 => x"ff4a4970",
   515 => x"c5c848d0",
   516 => x"7bd4c178",
   517 => x"7bbf976e",
   518 => x"80c1486e",
   519 => x"8dc17e70",
   520 => x"87f0ff05",
   521 => x"c448d0ff",
   522 => x"059a7278",
   523 => x"48c087c5",
   524 => x"c187e5c0",
   525 => x"e6f9c21e",
   526 => x"ecc4fe49",
   527 => x"7486c487",
   528 => x"c4fe059c",
   529 => x"48d0ff87",
   530 => x"c178c5c8",
   531 => x"7bc07bd3",
   532 => x"48c178c4",
   533 => x"48c087c2",
   534 => x"264d2626",
   535 => x"264b264c",
   536 => x"5b5e0e4f",
   537 => x"4b710e5c",
   538 => x"d80266cc",
   539 => x"f0c04c87",
   540 => x"87d8028c",
   541 => x"8ac14a74",
   542 => x"8a87d102",
   543 => x"8a87cd02",
   544 => x"d787c902",
   545 => x"fb497387",
   546 => x"87d087ea",
   547 => x"49c01e74",
   548 => x"7487dff9",
   549 => x"f949731e",
   550 => x"86c887d8",
   551 => x"0087fcfe",
   552 => x"c9e3c21e",
   553 => x"b9c149bf",
   554 => x"59cde3c2",
   555 => x"c348d4ff",
   556 => x"d0ff78ff",
   557 => x"78e1c848",
   558 => x"c148d4ff",
   559 => x"7131c478",
   560 => x"48d0ff78",
   561 => x"2678e0c0",
   562 => x"0000004f",
   563 => x"00000000",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
